* NGSPICE file created from housekeeping.ext - technology: gf180mcuC

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__fill_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__fill_2 VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__fillcap_4 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__fillcap_4 VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__fillcap_16 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__fillcap_16 VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__dffnsnq_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__dffnsnq_1 D SETN CLKN Q VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__fill_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__fill_1 VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__nor2_4 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__nor2_4 A1 A2 ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__dffsnq_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__dffsnq_1 D SETN CLK Q VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__aoi222_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__aoi222_1 A1 A2 B1 B2 C1 C2 ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__aoi22_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__aoi22_1 A1 A2 B1 B2 ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__nand4_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__nand4_1 A1 A2 A3 A4 ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__nand4_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__nand4_2 A1 A2 A3 A4 ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__fillcap_8 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__fillcap_8 VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__oai21_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__oai21_1 A1 A2 B ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__nor3_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__nor3_1 A1 A2 A3 ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__nand2_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__nand2_1 A1 A2 ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__dlyd_4 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__dlyd_4 I Z VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__and2_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__and2_1 A1 A2 Z VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__filltie abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__filltie VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__or2_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__or2_1 A1 A2 Z VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__nand2_4 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__nand2_4 A1 A2 ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__aoi21_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__aoi21_1 A1 A2 B ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__aoi211_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__aoi211_1 A1 A2 B C ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__nor2_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__nor2_1 A1 A2 ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__nor4_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__nor4_2 A1 A2 A3 A4 ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__dffq_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__dffq_1 D CLK Q VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 D RN CLK Q VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__nor2_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__nor2_2 A1 A2 ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__mux2_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__mux2_2 I0 I1 S Z VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__xor2_4 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__xor2_4 A1 A2 Z VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__oai31_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__oai31_2 A1 A2 A3 B ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__clkinv_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__clkinv_1 I ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__buf_8 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__buf_8 I Z VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__nand4_4 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__nand4_4 A1 A2 A3 A4 ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__or4_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__or4_2 A1 A2 A3 A4 Z VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__oai22_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__oai22_1 A1 A2 B1 B2 ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__and3_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__and3_1 A1 A2 A3 Z VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__dffsnq_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__dffsnq_2 D SETN CLK Q VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__nor4_4 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__nor4_4 A1 A2 A3 A4 ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__fillcap_32 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__fillcap_32 VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 I Z VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__endcap abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__endcap VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__nand3_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__nand3_1 A1 A2 A3 ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__dffrnq_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__dffrnq_2 D RN CLK Q VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__nor3_4 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__nor3_4 A1 A2 A3 ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__buf_12 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__buf_12 I Z VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 I Z VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__dffnrnq_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__dffnrnq_1 D RN CLKN Q VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__nand3_4 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__nand3_4 A1 A2 A3 ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__and4_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__and4_1 A1 A2 A3 A4 Z VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__aoi221_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__aoi221_1 A1 A2 B1 B2 C ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__oai32_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__oai32_1 A1 A2 A3 B1 B2 ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__oai21_4 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__oai21_4 A1 A2 B ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__inv_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__inv_1 I ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__oai21_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__oai21_2 A1 A2 B ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__nor4_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__nor4_1 A1 A2 A3 A4 ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__aoi222_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__aoi222_2 A1 A2 B1 B2 C1 C2 ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__oai211_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__oai211_1 A1 A2 B C ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__or2_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__or2_2 A1 A2 Z VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__nand2_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__nand2_2 A1 A2 ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__nor3_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__nor3_2 A1 A2 A3 ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__buf_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__buf_2 I Z VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__clkbuf_12 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__clkbuf_12 I Z VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__aoi211_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__aoi211_2 A1 A2 B C ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__aoi211_4 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__aoi211_4 A1 A2 B C ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__xor2_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__xor2_1 A1 A2 Z VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__aoi21_4 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__aoi21_4 A1 A2 B ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__oai31_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__oai31_1 A1 A2 A3 B ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__buf_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__buf_1 I Z VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__dffrnq_4 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__dffrnq_4 D RN CLK Q VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__or3_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__or3_1 A1 A2 A3 Z VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__clkinv_3 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__clkinv_3 I ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__or4_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__or4_1 A1 A2 A3 A4 Z VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__fillcap_64 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__fillcap_64 VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__inv_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__inv_2 I ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__or2_4 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__or2_4 A1 A2 Z VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__or3_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__or3_2 A1 A2 A3 Z VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__dffsnq_4 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__dffsnq_4 D SETN CLK Q VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__clkinv_12 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__clkinv_12 I ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__aoi221_4 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__aoi221_4 A1 A2 B1 B2 C ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__nand3_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__nand3_2 A1 A2 A3 ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__and2_4 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__and2_4 A1 A2 Z VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__aoi22_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__aoi22_2 A1 A2 B1 B2 ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__and4_4 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__and4_4 A1 A2 A3 A4 Z VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__mux2_4 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__mux2_4 I0 I1 S Z VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__or4_4 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__or4_4 A1 A2 A3 A4 Z VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__and3_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__and3_2 A1 A2 A3 Z VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__oai221_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__oai221_2 A1 A2 B1 B2 C ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__oai221_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__oai221_1 A1 A2 B1 B2 C ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__inv_3 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__inv_3 I ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__clkbuf_8 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__clkbuf_8 I Z VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__aoi21_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__aoi21_2 A1 A2 B ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__clkbuf_4 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__clkbuf_4 I Z VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__xnor2_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__xnor2_1 A1 A2 ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__oai22_4 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__oai22_4 A1 A2 B1 B2 ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 I Z VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__aoi221_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__aoi221_2 A1 A2 B1 B2 C ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__tieh abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__tieh Z VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__buf_16 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__buf_16 I Z VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__and2_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__and2_2 A1 A2 Z VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__buf_20 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__buf_20 I Z VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__oai211_4 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__oai211_4 A1 A2 B C ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__and4_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__and4_2 A1 A2 A3 A4 Z VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__clkinv_8 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__clkinv_8 I ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__inv_8 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__inv_8 I ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__oai33_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__oai33_1 A1 A2 A3 B1 B2 B3 ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__buf_3 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__buf_3 I Z VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__clkinv_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__clkinv_2 I ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__inv_4 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__inv_4 I ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__aoi22_4 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__aoi22_4 A1 A2 B1 B2 ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__oai32_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__oai32_2 A1 A2 A3 B1 B2 ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__aoi222_4 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__aoi222_4 A1 A2 B1 B2 C1 C2 ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__oai22_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__oai22_2 A1 A2 B1 B2 ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__xor2_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__xor2_2 A1 A2 Z VDD VSS
.ends

.subckt housekeeping VDD VSS debug_in debug_mode debug_oeb debug_out irq[0] irq[1]
+ irq[2] mask_rev_in[0] mask_rev_in[10] mask_rev_in[11] mask_rev_in[12] mask_rev_in[13]
+ mask_rev_in[14] mask_rev_in[15] mask_rev_in[16] mask_rev_in[17] mask_rev_in[18]
+ mask_rev_in[19] mask_rev_in[1] mask_rev_in[20] mask_rev_in[21] mask_rev_in[22] mask_rev_in[23]
+ mask_rev_in[24] mask_rev_in[25] mask_rev_in[26] mask_rev_in[27] mask_rev_in[28]
+ mask_rev_in[29] mask_rev_in[2] mask_rev_in[30] mask_rev_in[31] mask_rev_in[3] mask_rev_in[4]
+ mask_rev_in[5] mask_rev_in[6] mask_rev_in[7] mask_rev_in[8] mask_rev_in[9] mgmt_gpio_in[0]
+ mgmt_gpio_in[10] mgmt_gpio_in[11] mgmt_gpio_in[12] mgmt_gpio_in[13] mgmt_gpio_in[14]
+ mgmt_gpio_in[15] mgmt_gpio_in[16] mgmt_gpio_in[17] mgmt_gpio_in[18] mgmt_gpio_in[19]
+ mgmt_gpio_in[1] mgmt_gpio_in[20] mgmt_gpio_in[21] mgmt_gpio_in[22] mgmt_gpio_in[23]
+ mgmt_gpio_in[24] mgmt_gpio_in[25] mgmt_gpio_in[26] mgmt_gpio_in[27] mgmt_gpio_in[28]
+ mgmt_gpio_in[29] mgmt_gpio_in[2] mgmt_gpio_in[30] mgmt_gpio_in[31] mgmt_gpio_in[32]
+ mgmt_gpio_in[33] mgmt_gpio_in[34] mgmt_gpio_in[35] mgmt_gpio_in[36] mgmt_gpio_in[37]
+ mgmt_gpio_in[3] mgmt_gpio_in[4] mgmt_gpio_in[5] mgmt_gpio_in[6] mgmt_gpio_in[7]
+ mgmt_gpio_in[8] mgmt_gpio_in[9] mgmt_gpio_oeb[0] mgmt_gpio_oeb[10] mgmt_gpio_oeb[11]
+ mgmt_gpio_oeb[12] mgmt_gpio_oeb[13] mgmt_gpio_oeb[14] mgmt_gpio_oeb[15] mgmt_gpio_oeb[16]
+ mgmt_gpio_oeb[17] mgmt_gpio_oeb[18] mgmt_gpio_oeb[19] mgmt_gpio_oeb[1] mgmt_gpio_oeb[20]
+ mgmt_gpio_oeb[21] mgmt_gpio_oeb[22] mgmt_gpio_oeb[23] mgmt_gpio_oeb[24] mgmt_gpio_oeb[25]
+ mgmt_gpio_oeb[26] mgmt_gpio_oeb[27] mgmt_gpio_oeb[28] mgmt_gpio_oeb[29] mgmt_gpio_oeb[2]
+ mgmt_gpio_oeb[30] mgmt_gpio_oeb[31] mgmt_gpio_oeb[32] mgmt_gpio_oeb[33] mgmt_gpio_oeb[34]
+ mgmt_gpio_oeb[35] mgmt_gpio_oeb[36] mgmt_gpio_oeb[37] mgmt_gpio_oeb[3] mgmt_gpio_oeb[4]
+ mgmt_gpio_oeb[5] mgmt_gpio_oeb[6] mgmt_gpio_oeb[7] mgmt_gpio_oeb[8] mgmt_gpio_oeb[9]
+ mgmt_gpio_out[0] mgmt_gpio_out[10] mgmt_gpio_out[11] mgmt_gpio_out[12] mgmt_gpio_out[13]
+ mgmt_gpio_out[14] mgmt_gpio_out[15] mgmt_gpio_out[16] mgmt_gpio_out[17] mgmt_gpio_out[18]
+ mgmt_gpio_out[19] mgmt_gpio_out[1] mgmt_gpio_out[20] mgmt_gpio_out[21] mgmt_gpio_out[22]
+ mgmt_gpio_out[23] mgmt_gpio_out[24] mgmt_gpio_out[25] mgmt_gpio_out[26] mgmt_gpio_out[27]
+ mgmt_gpio_out[28] mgmt_gpio_out[29] mgmt_gpio_out[2] mgmt_gpio_out[30] mgmt_gpio_out[31]
+ mgmt_gpio_out[32] mgmt_gpio_out[33] mgmt_gpio_out[34] mgmt_gpio_out[35] mgmt_gpio_out[36]
+ mgmt_gpio_out[37] mgmt_gpio_out[3] mgmt_gpio_out[4] mgmt_gpio_out[5] mgmt_gpio_out[6]
+ mgmt_gpio_out[7] mgmt_gpio_out[8] mgmt_gpio_out[9] pad_flash_clk pad_flash_clk_oe
+ pad_flash_csb pad_flash_csb_oe pad_flash_io0_di pad_flash_io0_do pad_flash_io0_ie
+ pad_flash_io0_oe pad_flash_io1_di pad_flash_io1_do pad_flash_io1_ie pad_flash_io1_oe
+ pll90_sel[0] pll90_sel[1] pll90_sel[2] pll_bypass pll_dco_ena pll_div[0] pll_div[1]
+ pll_div[2] pll_div[3] pll_div[4] pll_ena pll_sel[0] pll_sel[1] pll_sel[2] pll_trim[0]
+ pll_trim[10] pll_trim[11] pll_trim[12] pll_trim[13] pll_trim[14] pll_trim[15] pll_trim[16]
+ pll_trim[17] pll_trim[18] pll_trim[19] pll_trim[1] pll_trim[20] pll_trim[21] pll_trim[22]
+ pll_trim[23] pll_trim[24] pll_trim[25] pll_trim[2] pll_trim[3] pll_trim[4] pll_trim[5]
+ pll_trim[6] pll_trim[7] pll_trim[8] pll_trim[9] porb pwr_ctrl_out qspi_enabled reset
+ ser_rx ser_tx serial_clock serial_data_1 serial_data_2 serial_load serial_resetn
+ spi_csb spi_enabled spi_sck spi_sdi spi_sdo spi_sdoenb spimemio_flash_clk spimemio_flash_csb
+ spimemio_flash_io0_di spimemio_flash_io0_do spimemio_flash_io0_oeb spimemio_flash_io1_di
+ spimemio_flash_io1_do spimemio_flash_io1_oeb spimemio_flash_io2_di spimemio_flash_io2_do
+ spimemio_flash_io2_oeb spimemio_flash_io3_di spimemio_flash_io3_do spimemio_flash_io3_oeb
+ trap uart_enabled user_clock wb_ack_o wb_adr_i[0] wb_adr_i[10] wb_adr_i[11] wb_adr_i[12]
+ wb_adr_i[13] wb_adr_i[14] wb_adr_i[15] wb_adr_i[16] wb_adr_i[17] wb_adr_i[18] wb_adr_i[19]
+ wb_adr_i[1] wb_adr_i[20] wb_adr_i[21] wb_adr_i[22] wb_adr_i[23] wb_adr_i[24] wb_adr_i[25]
+ wb_adr_i[26] wb_adr_i[27] wb_adr_i[28] wb_adr_i[29] wb_adr_i[2] wb_adr_i[30] wb_adr_i[31]
+ wb_adr_i[3] wb_adr_i[4] wb_adr_i[5] wb_adr_i[6] wb_adr_i[7] wb_adr_i[8] wb_adr_i[9]
+ wb_clk_i wb_cyc_i wb_dat_i[0] wb_dat_i[10] wb_dat_i[11] wb_dat_i[12] wb_dat_i[13]
+ wb_dat_i[14] wb_dat_i[15] wb_dat_i[16] wb_dat_i[17] wb_dat_i[18] wb_dat_i[19] wb_dat_i[1]
+ wb_dat_i[20] wb_dat_i[21] wb_dat_i[22] wb_dat_i[23] wb_dat_i[24] wb_dat_i[25] wb_dat_i[26]
+ wb_dat_i[27] wb_dat_i[28] wb_dat_i[29] wb_dat_i[2] wb_dat_i[30] wb_dat_i[31] wb_dat_i[3]
+ wb_dat_i[4] wb_dat_i[5] wb_dat_i[6] wb_dat_i[7] wb_dat_i[8] wb_dat_i[9] wb_dat_o[0]
+ wb_dat_o[10] wb_dat_o[11] wb_dat_o[12] wb_dat_o[13] wb_dat_o[14] wb_dat_o[15] wb_dat_o[16]
+ wb_dat_o[17] wb_dat_o[18] wb_dat_o[19] wb_dat_o[1] wb_dat_o[20] wb_dat_o[21] wb_dat_o[22]
+ wb_dat_o[23] wb_dat_o[24] wb_dat_o[25] wb_dat_o[26] wb_dat_o[27] wb_dat_o[28] wb_dat_o[29]
+ wb_dat_o[2] wb_dat_o[30] wb_dat_o[31] wb_dat_o[3] wb_dat_o[4] wb_dat_o[5] wb_dat_o[6]
+ wb_dat_o[7] wb_dat_o[8] wb_dat_o[9] wb_rstn_i wb_sel_i[0] wb_sel_i[1] wb_sel_i[2]
+ wb_sel_i[3] wb_stb_i wb_we_i
XFILLER_39_211 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_67_564 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_94_383 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_82_534 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_7963_ _7963_/D _7316_/Z _7977_/CLK _7963_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffnsnq_1
XFILLER_27_428 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_27_439 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_54_258 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6914_ _6955_/A4 _6935_/A2 _7202_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_4
X_7894_ _7894_/D _7901_/RN _7898_/CLK _7894_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffsnq_1
X_6845_ _7667_/Q _6885_/A2 _6647_/Z _7619_/Q _6887_/B1 _7683_/Q _6847_/A2 VDD VSS
+ gf180mcu_fd_sc_mcu7t5v0__aoi222_1
XFILLER_52_29 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_168_29 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3988_ _7625_/Q _5954_/A1 _6226_/A1 _7753_/Q _3989_/A4 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_6776_ _6776_/A1 _6776_/A2 _6776_/A3 _6776_/A4 _6777_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand4_1
XFILLER_164_801 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5727_ _5331_/Z _5727_/A2 _5437_/B _5619_/Z _5763_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand4_2
XFILLER_109_706 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_148_374 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_136_514 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_109_728 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_148_396 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5658_ _5669_/A1 _5179_/B _5658_/B _5674_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_5589_ _5589_/A1 _5589_/A2 _5589_/A3 _5590_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor3_1
XFILLER_2_505 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4609_ _4609_/A1 _7285_/A2 _4613_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_144_580 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_123_219 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_117_783 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
Xhold351 _7619_/Q hold351/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
X_7328_ _7901_/RN _4334_/Z _7328_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__and2_1
Xhold362 _7785_/Q hold362/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
Xhold340 _7642_/Q hold340/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
X_7259_ _7518_/Q _7259_/A2 _7261_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_132_753 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_104_444 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_89_144 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xhold373 _7769_/Q hold373/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
Xhold384 _7639_/Q hold384/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
Xhold395 _7362_/Q hold395/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
XFILLER_77_328 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_58_531 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_133_54 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_85_361 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_133_98 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_45_225 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_45_236 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_1800 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_61_707 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_165_2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1833 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1822 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1811 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_14_601 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1866 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1855 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1844 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_53_280 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1899 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1888 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1877 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_13_144 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_14_678 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_42_62 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_155_812 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_127_525 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_182_620 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_158_95 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_5_310 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_181_141 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_115_709 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_5_354 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_142_528 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_123_720 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_114_219 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_150_583 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_96_637 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_3_23 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_37_704 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_64_534 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_36_203 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_36_247 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4960_ _5797_/B _4965_/B _4960_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__or2_1
XFILLER_17_483 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_51_206 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3911_ _3911_/A1 _3911_/A2 _3911_/A3 _3911_/A4 _3917_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand4_1
X_4891_ hold607/Z _4892_/A2 _4892_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_177_425 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3842_ _3796_/Z hold113/Z hold114/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_4
XFILLER_60_784 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_20_615 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6630_ _7907_/Q _6633_/A2 _6664_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_4
XFILLER_80_2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6561_ _7902_/Q _7903_/Q _6561_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_164_108 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_146_812 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5512_ _5621_/B _5648_/B2 _5512_/B _5514_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_3773_ _4292_/B _3774_/A2 _7965_/Q _3774_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_6492_ _4460_/Z _6502_/A2 _6492_/B _7872_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_9_682 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_118_569 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5443_ _5621_/B _5648_/B2 _5629_/B _5572_/B _5444_/A4 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XFILLER_105_208 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5374_ _5405_/B _5504_/A3 _5577_/B2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_4325_ _4309_/S _4325_/A2 _4325_/B _7336_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_7113_ _7796_/Q _7190_/A2 _7190_/B1 _7618_/Q _7190_/C1 _7706_/Q _7116_/A2 VDD VSS
+ gf180mcu_fd_sc_mcu7t5v0__aoi222_1
XFILLER_113_296 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_86_136 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_7044_ _7623_/Q _7195_/B1 _7200_/B1 _7865_/Q _7048_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_4256_ _4256_/A1 _4256_/A2 _4256_/A3 _4256_/A4 _4263_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand4_1
XFILLER_67_361 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_47_29 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4187_ _4187_/A1 _4187_/A2 _4187_/A3 _4187_/A4 _4203_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor4_2
XFILLER_55_545 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_55_567 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7946_ _7946_/D _7949_/CLK _7946_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_1118 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1129 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1107 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_55_589 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7877_ _7877_/D _7901_/RN _7877_/CLK _7877_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_35_280 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_36_792 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6828_ _7927_/Q _7133_/S _6829_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_23_442 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_50_250 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_11_626 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_137_812 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_109_514 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6759_ _7728_/Q _6892_/B1 _6880_/B1 _7810_/Q _6766_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_128_21 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_109_525 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_163_141 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xhold170 _7438_/Q hold170/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
XFILLER_105_753 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
Xhold192 hold192/I _6225_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
Xhold181 _7655_/Q hold181/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
XFILLER_92_128 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_46_534 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2320 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_18_247 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_37_73 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2353 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2342 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2331 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_18_269 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2386 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2375 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2364 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1641 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1630 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2397 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_159_425 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1685 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1674 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1663 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1652 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1696 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_53_83 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_146_108 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_128_812 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_167_480 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_127_344 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_6_663 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_123_561 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_111_712 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5090_ _5692_/B _5285_/A3 _5424_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_2
XFILLER_123_594 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4110_ _4110_/I0 _7550_/Q _4427_/B _7550_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_4041_ _7719_/Q _6158_/A1 _4046_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_49_350 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_49_372 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_25_707 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_37_567 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7800_ _7800_/D _7901_/RN _7809_/CLK _7800_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffsnq_1
XFILLER_92_673 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5992_ _4454_/Z _6004_/A2 _5992_/B _7637_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_52_515 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_7731_ _7731_/D _7901_/RN _7755_/CLK _7731_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
X_4943_ _3728_/I _4900_/Z _4943_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__xor2_4
X_7662_ _7662_/D _7901_/RN _7797_/CLK _7662_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffsnq_1
XFILLER_32_250 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_33_762 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4874_ hold756/Z _4877_/A2 _4875_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_32_261 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6613_ _7915_/Q _6905_/A2 _6955_/A4 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_4
XFILLER_165_428 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_137_119 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_119_812 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7593_ _7593_/D input75/Z _7889_/CLK _8003_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
X_3825_ _4153_/A1 _4212_/A2 _6056_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_4
X_6544_ hold520/Z _6553_/A2 _6545_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_3756_ _4383_/A2 _3772_/S _4291_/A2 _3756_/B _3765_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai31_2
XFILLER_145_141 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6475_ _4460_/Z _6485_/A2 _6475_/B hold258/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_3687_ _7801_/Q _3687_/ZN VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_118_388 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5426_ _5712_/B _5534_/A2 _5691_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_1
Xoutput242 _7986_/Z mgmt_gpio_out[5] VDD VSS gf180mcu_fd_sc_mcu7t5v0__buf_8
Xoutput253 _4422_/I pad_flash_io0_oe VDD VSS gf180mcu_fd_sc_mcu7t5v0__buf_8
Xoutput220 _4404_/ZN mgmt_gpio_out[1] VDD VSS gf180mcu_fd_sc_mcu7t5v0__buf_8
Xoutput231 _7983_/Z mgmt_gpio_out[2] VDD VSS gf180mcu_fd_sc_mcu7t5v0__buf_8
X_5357_ _5357_/A1 _5643_/A2 _5667_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
Xoutput264 _7560_/Q pll_div[2] VDD VSS gf180mcu_fd_sc_mcu7t5v0__buf_8
Xoutput275 _7360_/Q pll_trim[13] VDD VSS gf180mcu_fd_sc_mcu7t5v0__buf_8
Xoutput286 _7354_/Q pll_trim[23] VDD VSS gf180mcu_fd_sc_mcu7t5v0__buf_8
XFILLER_181_18 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4308_ _3808_/Z _4308_/I1 _4308_/S _4308_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_101_211 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_99_283 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5288_ _5288_/A1 _5288_/A2 _5288_/A3 _5288_/A4 _5298_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand4_1
Xoutput297 _7572_/Q pwr_ctrl_out VDD VSS gf180mcu_fd_sc_mcu7t5v0__buf_8
X_7027_ _7027_/A1 _7210_/A2 _7027_/B _7433_/Q _7028_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi211_1
X_4239_ input20/Z _4239_/A2 _4774_/A1 _7474_/Q _4240_/A4 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_68_692 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_83_651 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_28_534 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_15_239 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_7929_ _7929_/D _7961_/RN _7940_/CLK _7929_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_169_712 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_130_66 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_90_37 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_70_389 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_11_423 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_24_795 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_51_570 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_128_108 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_128_2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_11_478 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_109_333 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_99_24 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_151_144 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_120_531 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_78_445 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_2_176 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_78_456 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_171_73 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_74_673 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_73_161 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_19_567 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_46_353 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2161 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2150 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_61_334 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_34_548 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2194 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2183 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2172 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1460 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_61_378 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_61_367 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1493 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1482 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1471 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_14_250 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_147_428 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4590_ hold661/Z _4593_/A2 _4591_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_30_776 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_174_247 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_127_141 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_142_100 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_6_460 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_182_291 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_142_122 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6260_ hold47/Z _6264_/A2 _6260_/B _7763_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_6191_ hold90/Z _6191_/A2 _6191_/B _7731_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_5211_ _3723_/I _4906_/S _5211_/A3 _4920_/Z _5373_/A4 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand4_4
XFILLER_43_2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5142_ _5309_/A1 _3723_/I _5006_/B _5254_/A2 _5545_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand4_4
XFILLER_142_199 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_130_339 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_69_445 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_69_423 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5073_ _4943_/Z _4993_/B _5663_/A1 _5077_/C VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor3_1
XFILLER_84_459 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4024_ _4024_/A1 _4024_/A2 _4024_/A3 _4024_/A4 _4025_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand4_1
XFILLER_80_621 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_5975_ _4454_/Z _5987_/A2 _5975_/B _7629_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_80_676 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4926_ _4926_/A1 _4926_/A2 _4926_/A3 _4926_/A4 _4926_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__or4_2
XFILLER_178_531 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7714_ _7714_/D _7901_/RN _7743_/CLK _7714_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_33_570 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_40_529 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_52_389 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4857_ _4454_/Z _4857_/A2 _4857_/B _7522_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_7645_ _7645_/D _7961_/RN _7645_/CLK _7645_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffsnq_1
XFILLER_176_29 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3808_ hold628/Z hold121/Z _7414_/Q _3808_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_60_29 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_7576_ _7576_/D _7961_/RN _7580_/CLK _7576_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
X_6527_ hold566/Z _6536_/A2 _6528_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_4788_ _7221_/A1 _4795_/S _4788_/B _7479_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_180_228 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_118_174 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3739_ _7344_/Q _3730_/Z _4383_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_6458_ _4460_/Z _6468_/A2 _6458_/B hold180/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_161_486 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_133_144 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6389_ hold265/Z _6400_/A2 hold266/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_121_306 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_5409_ _4993_/C _5099_/B _5645_/A3 _5409_/B2 _5411_/C VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai22_1
XFILLER_102_531 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_88_743 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_125_77 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_87_286 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_75_448 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_56_640 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_141_43 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_16_504 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_56_673 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_70_131 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_70_153 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_34_85 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_129_428 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_8_747 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_156_258 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_156_247 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_109_141 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_11_297 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_11_286 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_165_770 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_109_152 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_507 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_529 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_518 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_3_496 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_182_72 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_93_212 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_15_6 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_75_70 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_62_676 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5760_ _5617_/Z _5684_/Z _5760_/A3 _5760_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__and3_1
XFILLER_15_570 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_34_389 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4711_ _7442_/Q _4718_/A1 _4714_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_5691_ _5691_/A1 _5622_/Z _5691_/A3 _5691_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__and3_1
XTAP_1290 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_4642_ _3830_/Z hold47/Z _4643_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_7430_ hold70/Z _7901_/RN _7583_/CLK _7430_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_30_573 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_147_247 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
Xhold703 hold703/I _4509_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
X_7361_ _7361_/D _7961_/RN _7875_/CLK _7361_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffsnq_2
X_4573_ _4454_/Z _4573_/A2 _4573_/B _7392_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_7292_ _7901_/RN _4334_/Z _7292_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__and2_1
X_6312_ hold510/Z _6315_/A2 _6313_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
Xhold736 hold736/I _4456_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
Xhold714 _7403_/Q hold714/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
Xhold725 _7669_/Q hold725/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
XFILLER_170_261 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_170_250 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_115_144 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
Xhold747 _7604_/Q hold747/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
Xhold758 _7396_/Q hold758/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
X_6243_ _6243_/A1 _7285_/A2 _6247_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
Xhold769 _7732_/Q hold769/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
XFILLER_115_199 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_115_177 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_6174_ hold90/Z _6174_/A2 _6174_/B _7723_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_5125_ _5543_/C _5543_/B _5479_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_85_724 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_69_286 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5056_ _5199_/B _3727_/I _3728_/I _5369_/B _5087_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor4_4
XFILLER_111_383 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_38_640 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_57_459 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_84_267 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_4007_ hold124/Z hold25/Z _5817_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_4
XFILLER_55_29 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_52_120 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_80_484 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_80_473 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5958_ _4454_/Z _5970_/A2 _5958_/B _7621_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_4909_ _4925_/A1 _4923_/A1 _4914_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_166_534 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_5889_ hold577/Z _5902_/A2 _5890_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_21_551 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_7628_ _7628_/D _7901_/RN _7806_/CLK _7628_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffsnq_1
XFILLER_138_247 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_5_706 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_7559_ _7559_/D input75/Z _7567_/CLK _7559_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_106_144 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_161_283 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_121_114 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_106_188 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_422 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_136_98 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_96_69 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_96_58 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_76_702 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
Xhold41 hold41/I hold41/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
XFILLER_88_573 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
Xhold30 hold30/I hold30/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
XFILLER_75_212 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_488 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
Xhold74 hold74/I hold74/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
Xhold63 hold63/I hold63/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
XFILLER_152_64 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
Xhold52 hold52/I hold52/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
XFILLER_130_692 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xhold96 hold96/I hold96/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
Xhold85 hold85/I hold85/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
XFILLER_152_86 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_91_749 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_16_323 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_44_632 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
Xclkbuf_3_7__f_wb_clk_i clkbuf_0_wb_clk_i/Z _7958_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_45_73 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_44_676 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_71_495 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_16_389 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_351 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_340 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_12_540 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_362 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_157_567 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_12_584 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_145_729 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_6_34 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_152_250 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_99_805 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_112_103 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_140_489 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_120_191 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_54_407 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_81_215 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_19_172 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_35_621 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_47_470 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_6930_ _7914_/Q _7913_/Q _6599_/Z _6941_/A2 _7190_/B1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor4_4
Xclkbuf_leaf_6_csclk clkbuf_leaf_9_csclk/I _7895_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_23_805 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_34_120 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6861_ _7399_/Q _6894_/A2 _6891_/A2 _7407_/Q _6864_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_6792_ _7689_/Q _6884_/B1 _6792_/B _6792_/C _6800_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi211_1
X_5812_ _5812_/A1 _7285_/A2 _5816_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_35_676 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5743_ _5743_/A1 _5743_/A2 _5743_/A3 _5766_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_50_668 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_176_810 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_148_534 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5674_ _5674_/A1 _5674_/A2 _5674_/A3 _5773_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_30_392 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_4625_ _7991_/I _4652_/A1 _4628_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_129_770 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7413_ _7413_/D _7304_/Z _7977_/CLK _7413_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_2
XFILLER_144_740 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xhold500 _7866_/Q hold500/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
Xhold511 _7607_/Q hold511/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
X_4556_ _4448_/Z _4558_/A2 _4556_/B _7385_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_7344_ _7344_/D _7299_/Z _7977_/CLK _7344_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_2
Xhold522 _7891_/Q hold522/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
Xhold533 hold533/I _4519_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
Xhold544 hold544/I _4517_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
X_7275_ _7520_/Q _7275_/A2 _7275_/B1 _7519_/Q _7276_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_171_570 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_143_283 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_103_114 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_103_103 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
Xhold566 _7889_/Q hold566/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
Xhold577 _7999_/I hold577/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
Xhold555 _7358_/Q hold555/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
Xhold588 hold588/I _7495_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
XFILLER_1_219 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4487_ _4487_/A1 hold90/Z _4487_/B hold299/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_6226_ _6226_/A1 hold32/Z _6242_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_4
XFILLER_103_158 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xhold599 _7473_/Q hold599/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
X_6157_ hold90/Z _6157_/A2 _6157_/B _7715_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_106_68 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_860 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_871 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_5108_ _5661_/A1 _5797_/C _5647_/A2 _5672_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor3_4
XFILLER_85_554 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_58_768 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_882 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_893 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_57_212 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6088_ hold237/Z _6089_/A2 hold238/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_5039_ _5151_/A1 _5151_/A2 _5041_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_167_6 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_26_665 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_25_153 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_26_676 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_40_101 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_53_462 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_41_657 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_40_156 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_40_167 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_139_556 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_154_515 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_110_2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_134_250 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_150_721 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_135_795 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xinput120 wb_adr_i[3] _5006_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__buf_12
Xinput142 wb_dat_i[22] _7270_/B1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
Xinput131 wb_dat_i[12] _7260_/B1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
Xinput153 wb_dat_i[3] _7257_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_88_392 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xinput164 wb_sel_i[3] _7281_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_64_749 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_63_215 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_72_771 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_32_602 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_44_473 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_149_309 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_170 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_31_156 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XPHY_192 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_181 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_173_802 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_117_206 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_12_392 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_4410_ _7443_/Q user_clock _7584_/Q _4410_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_160_518 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5390_ _5660_/A2 _5390_/A2 _5701_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_126_751 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_172_389 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4341_ _7519_/Q _4438_/A2 _7514_/Q _4342_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_153_570 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_125_283 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_98_101 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_7060_ _7802_/Q _7191_/B1 _7190_/C1 _7704_/Q _7063_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_4272_ _7363_/Q _4505_/A1 _4569_/A1 _7391_/Q _4274_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_6011_ _4460_/Z _6021_/A2 _6011_/B hold30/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_86_318 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_67_543 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_67_532 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7962_ _7962_/D _7315_/Z _4031_/C2 hold11/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffnrnq_1
XFILLER_27_418 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_39_278 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_82_579 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_6913_ _7914_/Q _7913_/Q _6936_/A1 _6935_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand3_4
X_7893_ _7893_/D _7901_/RN _7893_/CLK _7893_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
X_6844_ _7805_/Q _6883_/A2 _6883_/B1 _7789_/Q _6884_/B1 _7691_/Q _6847_/A1 VDD VSS
+ gf180mcu_fd_sc_mcu7t5v0__aoi222_1
X_3987_ _7705_/Q _6124_/A1 _6107_/A1 _7697_/Q _3989_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_6775_ _7712_/Q _6885_/B1 _6890_/A2 _7640_/Q _6776_/A4 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_5726_ _5726_/A1 _5726_/A2 _5761_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_10_318 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_176_673 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_175_183 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5657_ _5706_/A1 _5657_/A2 _5657_/A3 _5657_/A4 _5657_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__and4_1
XFILLER_151_518 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_117_12 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5588_ _5673_/A2 _5566_/B _5588_/A3 _5733_/A3 _5589_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand4_1
X_4608_ _4454_/Z _4608_/A2 _4608_/B _7406_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_4539_ hold301/Z _4548_/A2 _4540_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_163_389 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_144_592 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_116_250 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xhold352 hold352/I _7619_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
Xhold330 _7784_/Q hold330/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
X_7327_ input75/Z _4334_/Z _7327_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__and2_1
Xhold341 hold341/I _7642_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
X_7258_ _7258_/A1 _7277_/B _7258_/B _7953_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi21_1
Xhold374 _7723_/Q hold374/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
XFILLER_104_434 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_89_123 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xhold363 _8001_/I hold363/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
Xhold385 hold385/I _7639_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
Xhold396 hold396/I _4504_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
XFILLER_104_467 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6209_ _6209_/A1 _7285_/A2 _6225_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_4
XFILLER_131_286 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_7189_ _7528_/Q _7189_/A2 _7189_/B1 _7522_/Q _7189_/C1 _7495_/Q _7192_/A1 VDD VSS
+ gf180mcu_fd_sc_mcu7t5v0__aoi222_1
XFILLER_133_66 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_133_33 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_690 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_100_673 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_39_790 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_45_215 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1834 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1823 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1812 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1801 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_159_618 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_158_2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1867 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1856 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1845 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_13_101 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1889 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1878 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_166_161 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_127_515 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_6_812 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_182_643 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_182_632 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_166_183 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_139_386 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_182_676 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_182_654 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_154_367 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_142_518 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_182_698 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_182_687 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_154_389 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_135_570 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_107_283 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_3_13 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_96_605 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_68_329 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_68_318 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_1_550 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_95_148 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_95_115 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_67_82 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_64_502 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_49_565 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
Xclkbuf_leaf_71_csclk _7961_/CLK _7650_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_37_738 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_91_354 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_83_70 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3910_ _7739_/Q _6192_/A1 _6107_/A1 _7699_/Q _3911_/A4 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_83_81 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xclkbuf_leaf_86_csclk _7396_/CLK _7756_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
X_4890_ _4448_/Z _4892_/A2 _4890_/B _7535_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_3841_ _4212_/A2 hold118/Z _6192_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_4
XFILLER_20_605 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_32_443 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_32_454 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3772_ input58/Z hold1/I _3772_/S _7966_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_6560_ _7902_/Q _6564_/B _6560_/B _7902_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_5511_ _5648_/A1 _5669_/B _5431_/B _5648_/B2 _5511_/C _5514_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi221_1
XFILLER_118_504 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_73_2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_157_183 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_157_161 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_145_312 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_118_526 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6491_ hold332/Z _6502_/A2 _6492_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_173_665 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_161_805 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5442_ _5319_/C _5563_/B2 _5687_/B _5319_/B _5692_/A2 _5629_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai32_1
X_5373_ _4906_/Z _5585_/A1 _5373_/A3 _5373_/A4 _5576_/B2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand4_2
XFILLER_99_421 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4324_ _7336_/Q _4309_/S _4325_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
Xclkbuf_leaf_24_csclk _7825_/CLK _7867_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_114_743 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_99_432 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7112_ _7682_/Q _7191_/A2 _7116_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_141_551 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_7043_ _7043_/A1 _7043_/A2 _7043_/A3 _7054_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_113_286 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_87_638 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4255_ _7748_/Q _6226_/A1 _6243_/A1 _7756_/Q _4256_/A4 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_1
Xclkbuf_leaf_39_csclk clkbuf_3_7__f_csclk/Z _7820_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
X_4186_ _4186_/A1 _4186_/A2 _4187_/A4 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_27_215 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_82_321 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_103_69 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7945_ _7945_/D _7949_/CLK _7945_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_1119 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1108 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_63_29 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_36_782 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_179_29 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7876_ _7876_/D _7961_/RN _7876_/CLK _7876_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
X_6827_ _7433_/Q _7926_/Q _6827_/B _6829_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_51_774 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_168_459 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_11_638 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_51_785 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6758_ _7794_/Q _6893_/A2 _6890_/B1 _7850_/Q _6766_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_6_108 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_164_621 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_5709_ _5709_/A1 _5709_/A2 _5710_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_6689_ _7791_/Q _6893_/A2 _6893_/B1 _7767_/Q _6692_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_12_33 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_164_676 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_164_687 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_128_88 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_128_66 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_117_570 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_88_37 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xhold171 hold171/I _7438_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
Xhold160 hold160/I _7706_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
Xhold193 hold193/I _7747_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
XFILLER_78_605 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
Xhold182 hold182/I _6030_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
XFILLER_144_98 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_92_118 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_86_682 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_58_384 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2310 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2343 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2332 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2321 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_33_207 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2387 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2376 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2354 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2365 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1642 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1631 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1620 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_33_229 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2398 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1675 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1664 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1653 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_774 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_53_40 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_169_51 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1697 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1686 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_53_73 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_169_73 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_155_621 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_139_161 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_154_120 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_143_805 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_182_484 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_154_164 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_154_153 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_5_141 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_5_152 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_123_551 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_150_392 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_123_584 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_69_638 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_110_234 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_96_479 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4040_ _7889_/Q _6520_/A1 hold108/I input64/Z _4052_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_64_321 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_92_685 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5991_ hold631/Z _6004_/A2 _5992_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_7730_ _7730_/D _7901_/RN _7753_/CLK _7730_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
X_4942_ _4920_/Z _4973_/A3 _4942_/B _5600_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_4
XFILLER_18_782 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_52_549 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_177_212 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7661_ _7661_/D _7901_/RN _7806_/CLK _7661_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffsnq_1
X_4873_ _4873_/A1 _7285_/A2 _4877_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_6612_ _6612_/I _7915_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_7592_ _7592_/D input75/Z _7592_/CLK _8002_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
X_3824_ hold19/Z _3787_/Z hold127/Z _3963_/A4 _4212_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand4_4
XFILLER_20_446 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_6543_ _4460_/Z _6553_/A2 _6543_/B hold188/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_3755_ _7413_/Q _3738_/Z _4291_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_145_120 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3686_ _7809_/Q _3686_/ZN VDD VSS gf180mcu_fd_sc_mcu7t5v0__inv_1
X_6474_ hold257/Z _6485_/A2 _6475_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_118_345 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_173_484 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_160_101 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_146_676 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_5425_ _5062_/Z _5176_/B _5425_/B _5437_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_2
Xoutput210 _4397_/Z mgmt_gpio_out[10] VDD VSS gf180mcu_fd_sc_mcu7t5v0__buf_8
XFILLER_160_112 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
Xoutput232 _8004_/Z mgmt_gpio_out[30] VDD VSS gf180mcu_fd_sc_mcu7t5v0__buf_8
Xoutput221 _7994_/Z mgmt_gpio_out[20] VDD VSS gf180mcu_fd_sc_mcu7t5v0__buf_8
Xoutput243 _4400_/Z mgmt_gpio_out[6] VDD VSS gf180mcu_fd_sc_mcu7t5v0__buf_8
X_5356_ _5094_/C _5356_/A2 _5356_/A3 _5356_/A4 _5359_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand4_1
Xoutput254 _8007_/Z pad_flash_io1_do VDD VSS gf180mcu_fd_sc_mcu7t5v0__buf_8
Xoutput276 _7361_/Q pll_trim[14] VDD VSS gf180mcu_fd_sc_mcu7t5v0__buf_8
XFILLER_0_807 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xoutput265 _7561_/Q pll_div[3] VDD VSS gf180mcu_fd_sc_mcu7t5v0__buf_8
X_4307_ _4306_/Z _7341_/Q _4309_/S _7341_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_141_381 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5287_ _5575_/A2 _5425_/B _5287_/B _5287_/C _5288_/A4 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XFILLER_101_223 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xoutput287 _7569_/Q pll_trim[24] VDD VSS gf180mcu_fd_sc_mcu7t5v0__buf_8
Xoutput298 _4215_/Z reset VDD VSS gf180mcu_fd_sc_mcu7t5v0__buf_8
XFILLER_102_757 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7026_ _7210_/A2 _7026_/A2 _7026_/A3 _7026_/A4 _7027_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor4_1
XFILLER_87_479 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4238_ _7920_/Q hold26/I _4238_/B1 input93/Z _4240_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_95_490 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_83_641 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4169_ _7847_/Q _6435_/A1 _4249_/A2 input15/Z _5881_/A1 _7587_/Q _4170_/A3 VDD VSS
+ gf180mcu_fd_sc_mcu7t5v0__aoi222_2
XFILLER_130_12 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_55_354 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_130_34 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_130_23 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_43_549 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7928_ _7928_/D _7961_/RN _7938_/CLK _7928_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_55_398 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_23_240 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_168_212 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7859_ _7859_/D _7901_/RN _7900_/CLK _7859_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_169_779 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_139_43 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_137_621 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_109_323 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_7_428 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_139_65 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_23_98 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_136_153 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_152_646 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_3_2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_132_370 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_105_584 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_132_392 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_171_63 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_93_438 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_47_811 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_19_557 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_46_321 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_69 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2162 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2151 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2140 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_34_538 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2195 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2184 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2173 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1450 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_61_357 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_15_763 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_159_212 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1483 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1472 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1461 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_9_34 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_42_560 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1494 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_9_78 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_30_744 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_128_676 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5210_ _5087_/C _4914_/Z _5210_/A3 _5210_/B _5373_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai31_2
XFILLER_155_495 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_143_657 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6190_ hold195/Z _6191_/A2 _6191_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_130_318 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5141_ _3722_/I _5087_/C _5394_/A1 _5006_/C _5176_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor4_4
XFILLER_130_329 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_36_2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5072_ _5476_/B _5689_/A1 _5072_/B _5072_/C _5106_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_111_554 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_69_468 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4023_ _7810_/Q _6350_/A1 _6226_/A1 _7752_/Q _4024_/A4 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_56_129 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_65_641 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_37_354 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_37_398 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7713_ _7713_/D _7901_/RN _7753_/CLK _7713_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
X_5974_ hold693/Z _5987_/A2 _5975_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_4925_ _4925_/A1 input96/Z _4926_/A4 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_100_37 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4856_ hold590/Z _4857_/A2 _4857_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_7644_ _7644_/D _7961_/RN _7648_/CLK _7644_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffsnq_1
XFILLER_165_215 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_159_790 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_3807_ _7340_/Q _4383_/A1 _4308_/I1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_21_799 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_7575_ _7575_/D _7961_/RN _7580_/CLK _7575_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_165_248 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_119_654 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6526_ _4460_/Z _6536_/A2 _6526_/B hold190/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_4787_ _7479_/Q _4795_/S _4788_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_174_771 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_134_602 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3738_ _7344_/Q _3730_/Z _3738_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__and2_1
X_3669_ hold28/I _7253_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_118_186 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6457_ hold178/Z _6468_/A2 hold179/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_5408_ _5585_/A1 _5608_/B _5621_/B _5759_/A1 _5408_/C _5413_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi221_1
X_6388_ _4454_/Z _6400_/A2 _6388_/B _7823_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_5339_ _5200_/B _3727_/I _4915_/Z _5433_/C _5618_/B1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand4_4
XFILLER_114_392 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_659 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_125_89 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_48_619 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7009_ _7848_/Q _7193_/A2 _7193_/C1 _7726_/Q _7193_/B1 _7630_/Q _7016_/A1 VDD VSS
+ gf180mcu_fd_sc_mcu7t5v0__aoi222_1
XFILLER_18_43 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_28_321 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
Xclkbuf_3_6__f_wb_clk_i clkbuf_0_wb_clk_i/Z _4411_/I1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_141_77 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_83_471 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_71_633 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_16_527 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_28_387 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_141_99 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_71_655 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_43_357 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_70_176 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_34_53 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_140_2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_11_221 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_51_390 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_109_131 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_125_613 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_180_763 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_140_605 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_112_318 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_519 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_508 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_182_95 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_120_351 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_94_747 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_93_224 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_59_490 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_47_641 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_19_343 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_19_365 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_46_140 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_47_674 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_74_471 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_62_633 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_61_132 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_4710_ _4718_/A1 hold58/Z _4710_/B hold59/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_5690_ _5690_/A1 _5757_/A2 _5691_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_91_70 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1291 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1280 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_4641_ _7995_/I _4652_/A1 _4644_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_147_215 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_128_451 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_116_602 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7360_ _7360_/D _7961_/RN _7370_/CLK _7360_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffsnq_2
X_4572_ hold591/Z _4573_/A2 _4573_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_143_432 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7291_ _7901_/RN _4334_/Z _7291_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_115_112 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6311_ hold47/Z _6315_/A2 _6311_/B _7787_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
Xhold737 hold737/I _7348_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
Xhold726 _7556_/Q hold726/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
Xhold704 hold704/I _7364_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
Xhold715 _7405_/Q hold715/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
X_6242_ hold90/Z _6242_/A2 _6242_/B _7755_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_171_785 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xhold759 _7716_/Q hold759/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
XFILLER_115_156 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
Xhold748 _7758_/Q hold748/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
XFILLER_131_638 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_131_627 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6173_ hold374/Z _6174_/A2 _6174_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_69_221 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5124_ _5533_/A1 _5543_/B _5540_/B1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_97_585 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5055_ _3728_/I _5369_/B _5421_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_4
X_4006_ _7858_/Q _6452_/A1 _4035_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_93_780 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_1_90 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_53_622 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_25_346 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_25_357 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_111_58 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_80_463 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5957_ hold649/Z _5970_/A2 _5958_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_52_176 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4908_ _5302_/A1 _4365_/Z _5015_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__or2_2
XFILLER_139_716 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_40_327 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5888_ _4448_/Z _5902_/A2 _5888_/B _7588_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_7627_ _7627_/D _7961_/RN _7627_/CLK _7627_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
X_4839_ _5678_/A1 _7280_/A2 _7279_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_2
XFILLER_181_505 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7558_ _7558_/D input75/Z _7558_/CLK _7558_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_4_206 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_119_495 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6509_ _4460_/Z _6519_/A2 _6509_/B _7880_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_20_33 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7489_ _7489_/D _7912_/CLK _7489_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_136_33 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_136_44 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_122_605 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_136_77 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_96_37 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xhold31 hold31/I hold31/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
XFILLER_88_585 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
Xhold20 hold20/I hold20/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
XFILLER_29_42 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
Xhold42 hold42/I hold42/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
Xhold64 hold64/I hold64/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
XFILLER_88_596 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_76_747 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xhold75 hold75/I hold75/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
Xhold97 hold97/I hold97/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
Xhold86 hold86/I hold86/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
XFILLER_28_140 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_29_641 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_28_195 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_43_132 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_352 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_341 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_330 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_363 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_169_373 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_129_215 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_129_204 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_61_73 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_61_62 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_8_534 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_177_73 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_157_579 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_8_589 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_153_730 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_125_421 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_113_638 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_3_283 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_94_511 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_79_563 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_94_522 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_94_544 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_94_566 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_82_717 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_75_780 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_34_132 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_6860_ _7476_/Q _6880_/C2 _6892_/A2 _7385_/Q _6860_/C _6873_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi221_1
XFILLER_47_493 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6791_ _6791_/A1 _6791_/A2 _6791_/A3 _6792_/C VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_62_463 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_22_316 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5811_ _4454_/Z _5811_/A2 _5811_/B _7547_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_5742_ _5742_/A1 _5506_/C _5550_/C _5742_/A4 _5743_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor4_1
XFILLER_22_327 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_34_187 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_50_658 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5673_ _5673_/A1 _5673_/A2 _5673_/A3 _5673_/A4 _5754_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand4_2
XFILLER_175_354 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4624_ _4652_/A1 hold101/Z _4624_/B hold102/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_7412_ _7412_/D _7303_/Z _7977_/CLK _7412_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_144_730 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7343_ _7343_/D _7298_/Z _4031_/C2 _7343_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
Xhold501 _7778_/Q hold501/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
X_4555_ hold719/Z _4558_/A2 _4556_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_104_605 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xhold523 _7835_/Q hold523/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
Xhold534 hold534/I _7369_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
Xhold545 hold545/I _7368_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
Xhold512 _7649_/Q hold512/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
X_7274_ _7518_/Q _7274_/A2 _7276_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
Xhold567 _7749_/Q hold567/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
X_4486_ hold90/Z _4753_/I1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_116_498 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_104_638 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xhold556 hold556/I _4496_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
Xhold578 _7388_/Q hold578/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
X_6225_ hold90/Z _6225_/A2 _6225_/B hold193/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_106_14 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_103_137 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xhold589 _7895_/Q hold589/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
X_6156_ hold204/Z _6157_/A2 _6157_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_106_58 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_97_371 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_850 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_861 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_5107_ _5319_/C _5692_/B _5563_/B2 _5591_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor3_2
XFILLER_66_29 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_58_747 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_872 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_883 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_894 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_6087_ hold68/Z _6089_/A2 _6087_/B _7682_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_111_192 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_85_566 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5038_ _5038_/A1 _5038_/A2 _5038_/A3 _5106_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_38_460 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_122_68 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_14_806 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_81_783 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_53_485 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_6989_ _7895_/Q _7197_/A2 _6938_/I _7855_/Q _6990_/A4 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_40_124 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_178_170 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_166_321 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_21_371 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_40_179 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_182_803 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_147_43 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_181_357 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_103_2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_31_87 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_147_98 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_150_744 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xinput110 wb_adr_i[23] _5224_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__buf_2
Xinput143 wb_dat_i[23] _7274_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
Xinput132 wb_dat_i[13] _7265_/B1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
Xinput154 wb_dat_i[4] _7262_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
Xinput121 wb_adr_i[4] _3728_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_12
XFILLER_0_286 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_102_192 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
Xinput165 wb_stb_i _4366_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_48_246 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_44_463 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_72_61 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_16_176 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_31_124 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XPHY_160 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_32_669 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_193 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_182 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_171 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_172_302 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_157_354 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_157_398 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_8_386 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_172_346 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_126_763 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_99_603 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4340_ _4340_/I _7518_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_141_700 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_140_210 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_98_124 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4271_ _4271_/A1 _4271_/A2 _4271_/A3 _4281_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_98_179 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6010_ _7646_/Q _6021_/A2 _6011_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_100_129 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_94_396 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_82_525 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_7961_ _7961_/D _7961_/RN _7961_/CLK _7961_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
X_7892_ _7892_/D _7901_/RN _7893_/CLK _7892_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
X_6912_ _6953_/A1 _6950_/A1 _6955_/A4 _7200_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor3_4
X_6843_ _6843_/A1 _6843_/A2 _6843_/A3 _6848_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_63_783 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_23_647 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_35_485 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_35_496 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_149_800 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3986_ _7721_/Q _6158_/A1 _6248_/A1 _7763_/Q _3989_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_6774_ _7720_/Q _6881_/A2 _6881_/B1 _7696_/Q _6776_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_50_455 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_148_321 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5725_ _5725_/A1 _5725_/A2 _5725_/A3 _5726_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_22_179 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_176_663 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_136_516 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5656_ _5656_/A1 _5656_/A2 _5748_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_148_387 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4607_ hold610/Z _4608_/A2 _4608_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_163_357 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xhold320 _7810_/Q hold320/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
X_5587_ _5062_/Z _5425_/B _5587_/B _5587_/C _5733_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi211_2
XFILLER_117_763 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_4538_ _4460_/Z _4548_/A2 _4538_/B hold115/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
Xhold331 _7727_/Q hold331/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
XFILLER_117_24 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xhold353 _7699_/Q hold353/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
Xhold342 _7611_/Q hold342/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
X_7326_ input75/Z _4334_/Z _7326_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__and2_1
X_7257_ _7257_/A1 _7280_/A2 _7277_/B _7257_/C _7258_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi211_1
X_4469_ _7969_/Q _7506_/Q hold40/Z hold41/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_4
Xhold375 _7765_/Q hold375/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
Xhold386 _7770_/Q hold386/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
Xhold364 _7865_/Q hold364/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
X_6208_ hold90/Z _6208_/A2 _6208_/B _7739_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
Xhold397 hold397/I _7362_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
X_7188_ _7757_/Q _7188_/A2 _7198_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_6139_ hold354/Z _6140_/A2 _6140_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_680 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_691 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_73_503 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_39_780 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_45_227 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_61_709 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1824 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1813 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1802 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_26_463 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1857 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1846 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1835 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_81_580 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_53_260 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1879 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1868 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_167_641 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_13_168 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_41_499 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_139_365 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_139_354 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_139_343 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_158_75 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_142_508 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_123_722 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_150_530 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
Xclkbuf_leaf_5_csclk clkbuf_leaf_9_csclk/I _7887_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_96_628 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_1_540 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_110_427 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_89_691 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_49_533 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_92_812 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_76_363 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_64_558 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_45_783 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_17_496 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_149_118 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3840_ _3801_/Z hold117/Z hold24/Z hold274/I hold118/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand4_4
X_3771_ hold1/I hold5/I _3772_/S _7967_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_32_488 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_157_140 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5510_ _5621_/B _5510_/A2 _5510_/B _5752_/C _5514_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XFILLER_173_611 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_172_110 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_157_173 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6490_ _4454_/Z _6502_/A2 _6490_/B _7871_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_5441_ _5591_/A2 _5501_/A2 _5613_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_145_357 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_66_2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5372_ _5375_/A4 _5382_/A3 _5372_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__or2_1
XFILLER_172_176 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4323_ input58/Z _4383_/A1 _4323_/B _4325_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_7111_ _7111_/I _7115_/C VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_86_105 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7042_ _7897_/Q _7197_/A2 _7195_/C1 _7873_/Q _7043_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_99_499 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4254_ _7846_/Q _6435_/A1 _4609_/A1 _7407_/Q _4256_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_95_661 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4185_ _7879_/Q _6503_/A1 _6486_/A1 _7871_/Q _6124_/A1 _7701_/Q _4186_/A2 VDD VSS
+ gf180mcu_fd_sc_mcu7t5v0__aoi222_1
XFILLER_83_812 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_28_739 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_7944_ _7944_/D _7944_/CLK _7944_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_43_709 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1109 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_63_591 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7875_ _7875_/D _7961_/RN _7875_/CLK _7875_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
X_6826_ _6826_/A1 _6767_/C _6826_/B _7433_/Q _6827_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XFILLER_23_444 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_168_449 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_149_641 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6757_ _7133_/S _6757_/A2 _6757_/B _7924_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_10_105 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_23_499 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5708_ _5104_/B _5708_/A2 _5708_/B _5710_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_3969_ _7891_/Q _6520_/A1 _5920_/A1 _7609_/Q _3981_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_148_162 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_6688_ _7775_/Q _6891_/C1 _6692_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_148_195 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_5639_ _5656_/A1 _5639_/A2 _5639_/B _5639_/C _5640_/B2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XFILLER_128_34 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_124_508 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_12_67 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_132_530 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
Xhold161 _7597_/Q hold161/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
Xhold150 hold150/I _7606_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
XFILLER_2_348 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7309_ input75/Z _4334_/Z _7309_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__and2_1
Xhold194 _7755_/Q hold194/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
Xhold172 _7600_/Q hold172/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
XFILLER_105_777 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xhold183 hold183/I _7655_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
XFILLER_120_747 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_92_108 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_74_812 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_37_42 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_46_503 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2311 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2300 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_170_2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_85_171 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_18_238 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2344 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2333 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2322 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_37_86 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_46_569 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2377 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2355 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2366 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1632 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1621 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1610 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_61_539 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_14_400 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_27_783 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2399 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2388 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1676 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1665 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1654 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1643 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_41_241 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1687 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1698 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_53_96 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_174_408 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_155_611 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_182_452 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_182_441 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_182_430 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_127_357 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_154_176 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_127_368 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_108_560 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_6_676 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_123_541 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_68_105 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_110_246 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_96_458 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_84_609 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_65_812 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_37_514 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_94_81 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_91_141 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5990_ _4448_/Z _6004_/A2 _5990_/B _7636_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_25_709 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4941_ _5210_/A3 _4974_/A3 _4941_/B _4941_/C _4951_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi211_4
XFILLER_64_399 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7660_ _7660_/D _7901_/RN _7852_/CLK _7660_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffsnq_1
X_4872_ _4454_/Z _4872_/A2 _4872_/B _7528_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_33_753 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_178_747 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_3823_ _3817_/I _4153_/A1 _6039_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_4
XFILLER_32_252 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6611_ _7915_/Q _6611_/A2 _6611_/B _6612_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_7591_ _7591_/D input75/Z _7865_/CLK _8001_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_20_458 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_158_460 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6542_ hold187/Z _6553_/A2 _6543_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_3754_ _7975_/Q _7974_/Q _4291_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_2
X_3685_ _7817_/Q _3685_/ZN VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_6473_ _4454_/Z _6485_/A2 _6473_/B _7863_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
Xoutput200 _4391_/ZN mgmt_gpio_oeb[36] VDD VSS gf180mcu_fd_sc_mcu7t5v0__buf_8
X_5424_ _5424_/A1 _5575_/A2 _5424_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_173_496 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xoutput233 _8005_/Z mgmt_gpio_out[31] VDD VSS gf180mcu_fd_sc_mcu7t5v0__buf_8
Xoutput211 _7988_/Z mgmt_gpio_out[11] VDD VSS gf180mcu_fd_sc_mcu7t5v0__buf_8
Xoutput222 _7995_/Z mgmt_gpio_out[21] VDD VSS gf180mcu_fd_sc_mcu7t5v0__buf_8
Xoutput244 _7987_/Z mgmt_gpio_out[7] VDD VSS gf180mcu_fd_sc_mcu7t5v0__buf_8
X_5355_ _5680_/A1 _5768_/A3 _5546_/B1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
Xoutput255 _4420_/I pad_flash_io1_ie VDD VSS gf180mcu_fd_sc_mcu7t5v0__buf_8
Xoutput266 _7562_/Q pll_div[4] VDD VSS gf180mcu_fd_sc_mcu7t5v0__buf_8
Xoutput277 _7362_/Q pll_trim[15] VDD VSS gf180mcu_fd_sc_mcu7t5v0__buf_8
XFILLER_160_179 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_4306_ _4306_/A1 _4306_/A2 _4306_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_5286_ _4996_/Z _5424_/A1 _5733_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_102_747 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_87_425 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xoutput288 _7570_/Q pll_trim[25] VDD VSS gf180mcu_fd_sc_mcu7t5v0__buf_8
Xoutput299 _4429_/Z ser_rx VDD VSS gf180mcu_fd_sc_mcu7t5v0__buf_8
X_7025_ _7025_/A1 _7025_/A2 _7025_/A3 _7025_/A4 _7026_/A4 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand4_1
XFILLER_101_235 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_87_447 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4237_ _7684_/Q _6090_/A1 _5874_/A1 _7585_/Q _4240_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_74_108 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_68_672 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_56_812 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xclkbuf_3_5__f_wb_clk_i clkbuf_0_wb_clk_i/Z _7545_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_74_29 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_28_536 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4168_ _7613_/Q _5937_/A1 _4831_/A1 _7505_/Q _4848_/A1 _7510_/Q _4170_/A2 VDD VSS
+ gf180mcu_fd_sc_mcu7t5v0__aoi222_2
X_4099_ _7776_/Q _6282_/A1 _6469_/A1 _7864_/Q _4100_/A4 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_82_141 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_70_303 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_55_366 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7927_ _7927_/D _7961_/RN _7949_/CLK _7927_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_169_725 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_90_17 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7858_ _7858_/D _7901_/RN _7898_/CLK _7858_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_70_369 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_70_358 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_24_742 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_142_6 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6809_ _7844_/Q _6894_/A2 _6891_/A2 _7828_/Q _6812_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_7789_ _7789_/D _7901_/RN _7900_/CLK _7789_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_11_425 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_177_780 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_139_55 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_137_611 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_11_469 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_149_493 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_128_4 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_109_357 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xclkbuf_leaf_70_csclk _7961_/CLK _7648_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_164_463 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_151_135 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_151_124 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_2_112 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_132_382 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_120_500 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_105_574 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xclkbuf_leaf_85_csclk _7396_/CLK _7874_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_93_428 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_171_86 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_101_780 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_19_547 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_104_80 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_73_141 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_37 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2152 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2141 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2130 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2185 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2174 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2163 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1451 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1440 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_15_753 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2196 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_159_224 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1484 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1473 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1462 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_14_263 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_42_572 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1495 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_175_728 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
Xclkbuf_leaf_38_csclk clkbuf_3_7__f_csclk/Z _7812_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_170_400 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_182_282 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_127_198 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_89_70 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5140_ _5543_/C _5498_/A2 _5498_/B _5187_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor3_1
XFILLER_142_179 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_123_371 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_123_382 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_97_712 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_96_211 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_69_425 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5071_ _5608_/A1 _5608_/B _5475_/B _5066_/Z _5071_/C _5072_/C VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi221_1
XFILLER_29_2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_111_566 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4022_ input39/Z _5903_/A1 _6316_/A1 _7794_/Q _4024_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_38_812 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_56_108 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_84_439 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_37_333 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5973_ _4448_/Z _5987_/A2 _5973_/B _7628_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_64_185 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_4924_ _4924_/A1 _4924_/A2 _4924_/A3 _4924_/A4 _4926_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand4_1
X_7712_ _7712_/D _7901_/RN _7812_/CLK _7712_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_80_678 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_40_509 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_100_16 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_21_712 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4855_ _4448_/Z _4857_/A2 _4855_/B _7521_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_20_233 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7643_ _7643_/D _7961_/RN _7643_/CLK _7643_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
X_3806_ _3801_/S hold754/Z _3806_/B _3864_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi21_4
XFILLER_119_600 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7574_ hold13/Z _7901_/RN _7802_/CLK _7982_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
X_4786_ _7219_/A1 _4795_/S _4786_/B _7478_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_181_709 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6525_ hold189/Z _6536_/A2 _6526_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_3737_ _7346_/Q _7344_/Q _3774_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_146_463 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_106_305 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3668_ hold34/I _7248_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_161_411 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_119_699 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_118_198 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_118_176 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_109_58 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_106_316 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6456_ _4454_/Z _6468_/A2 _6456_/B _7855_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_69_29 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5407_ _5782_/A1 _5407_/A2 _5407_/A3 _5414_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_133_168 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6387_ hold667/Z _6400_/A2 _6388_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_161_499 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5338_ _5338_/A1 _5421_/B1 _5779_/B1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_114_371 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_85_17 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_102_566 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5269_ _5624_/A1 _5624_/B _5586_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_7008_ _7008_/A1 _7008_/A2 _7008_/A3 _7008_/A4 _7026_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand4_1
XFILLER_87_288 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_75_428 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_29_812 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_18_33 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_55_141 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_71_645 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_24_594 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_133_2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_149_290 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_11_288 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_7_215 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_171_219 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_165_783 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_166_64 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_164_282 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_137_496 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_124_124 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_109_198 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_166_86 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_124_135 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_124_179 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_79_712 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_509 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_3_487 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_105_382 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_59_73 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_94_737 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_38_108 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_120_396 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_93_236 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_78_299 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_75_50 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_46_174 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_61_144 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_148_717 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_1292 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1281 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1270 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_30_531 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4640_ _4652_/A1 hold64/Z _4640_/B hold65/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_175_558 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_163_709 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_30_575 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_128_463 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6310_ hold521/Z _6315_/A2 _6311_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_4571_ _4448_/Z _4573_/A2 _4571_/B _7391_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
Xhold727 hold727/I _7556_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
Xhold705 _7557_/Q hold705/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
Xhold716 _7563_/Q hold716/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
X_7290_ input75/Z _4334_/Z _7290_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__and2_1
X_6241_ hold194/Z _6242_/A2 _6242_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
Xhold738 _7894_/Q hold738/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
Xhold749 _7525_/Q hold749/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
XFILLER_170_263 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_143_499 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6172_ hold68/Z _6174_/A2 _6172_/B _7722_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_115_168 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5123_ _4953_/Z _5139_/A1 _5014_/Z _5543_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand3_4
XFILLER_97_531 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5054_ _5199_/B _3727_/I _5054_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__or2_2
XFILLER_57_428 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_84_247 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4005_ _7882_/Q _6503_/A1 _6005_/A1 _7648_/Q _4024_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_93_792 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_52_122 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5956_ _4448_/Z _5970_/A2 _5956_/B _7620_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_4907_ _5302_/A1 _5224_/A3 _5224_/A4 _5016_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor3_4
X_5887_ hold665/Z _5902_/A2 _5888_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_52_188 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_4838_ _7516_/Q _5301_/B _5520_/C VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_4
XFILLER_166_525 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_7626_ _7626_/D _7961_/RN _7643_/CLK _7626_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_153_219 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7557_ _7557_/D input75/Z _7565_/CLK _7557_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffsnq_1
X_4769_ _4769_/A1 _7285_/A2 _4773_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_174_591 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_147_783 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_146_282 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_106_124 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_6508_ hold326/Z _6519_/A2 _6509_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_7488_ _7488_/D _7912_/CLK _7488_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_162_764 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_161_230 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_6439_ _4454_/Z _6451_/A2 _6439_/B _7847_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_136_56 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_106_179 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_102_330 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_88_531 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_88_520 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
Xhold10 hold10/I hold10/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
Xhold32 hold32/I hold32/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
XFILLER_88_575 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_457 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_29_32 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
Xhold21 hold21/I hold21/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
XFILLER_48_417 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
Xhold43 hold43/I hold43/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
Xhold65 hold65/I hold65/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
XFILLER_152_33 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_29_65 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xhold98 hold98/I hold98/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
Xhold76 hold76/I hold76/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
Xhold87 hold87/I hold87/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
XFILLER_16_347 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_43_144 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_342 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_331 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_320 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_101_70 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_364 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_353 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_12_531 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_177_30 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_125_411 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_4_741 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_125_499 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_125_477 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_112_105 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_112_149 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_106_680 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_140_469 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_94_534 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_39_428 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_19_141 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_75_770 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_62_431 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_62_420 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_35_634 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6790_ _7753_/Q _6644_/Z _6885_/B1 _7713_/Q _6791_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_62_475 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5810_ hold611/Z _5811_/A2 _5811_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_5741_ _5741_/A1 _4993_/B _5741_/A3 _5741_/B _5742_/A4 VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai31_1
XFILLER_96_2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_176_812 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_175_311 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5672_ _5179_/B _5672_/A2 _5793_/A2 _5606_/B _5673_/A4 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_7411_ _7411_/D _7302_/Z _7977_/CLK _7411_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffsnq_2
XFILLER_175_377 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4623_ hold100/Z _3830_/Z _4623_/B hold101/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_7342_ _7342_/D _7297_/Z _4031_/C2 _7342_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
Xhold502 _7793_/Q hold502/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
XFILLER_129_783 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_128_282 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4554_ _4554_/A1 _7285_/A2 _4558_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_7273_ _7273_/A1 _7277_/B _7273_/B _7956_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi21_1
Xhold524 _7883_/Q hold524/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
XFILLER_7_590 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
Xhold535 _7361_/Q hold535/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
Xhold513 hold513/I _7649_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
Xhold568 _7725_/Q hold568/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
X_4485_ _7972_/Q _7506_/Q hold89/Z hold90/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_4
X_6224_ hold191/Z _6225_/A2 hold192/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_131_414 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
Xhold546 _7615_/Q hold546/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
Xhold557 hold557/I _7358_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
Xhold579 _7471_/Q hold579/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
XFILLER_131_458 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_131_425 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6155_ hold68/Z _6157_/A2 _6155_/B _7714_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_106_37 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_100_812 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_97_361 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_840 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_851 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_862 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_6086_ hold408/Z _6089_/A2 _6087_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_5106_ _5106_/A1 _5106_/A2 _5106_/A3 _5106_/A4 _5115_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor4_1
XTAP_873 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_884 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_895 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_5037_ _5585_/A1 _5658_/B _5608_/B _5669_/A1 _5037_/C _5038_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi221_1
XFILLER_85_578 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_85_556 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_122_47 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_26_623 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_80_250 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_25_144 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_15_34 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_41_637 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6988_ _7887_/Q _7196_/A2 _7196_/B1 _7637_/Q _6990_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_167_812 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5939_ _4448_/Z _5953_/A2 _5939_/B _7612_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_40_136 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_40_158 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_127_709 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7609_ _7609_/D _7961_/RN _7694_/CLK _7609_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_31_77 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_162_550 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_134_252 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_150_756 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_107_499 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xinput111 wb_adr_i[24] _4370_/A4 VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
Xinput100 wb_adr_i[14] _4922_/A4 VDD VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_122_458 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_76_501 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xinput144 wb_dat_i[24] _7240_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
Xinput133 wb_dat_i[14] _7269_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
Xinput122 wb_adr_i[5] _5369_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__buf_12
XFILLER_163_98 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_76_534 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
Xinput166 wb_we_i _3658_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
Xinput155 wb_dat_i[5] _7267_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_76_567 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_17_623 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_44_431 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_56_291 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_44_442 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_112_91 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_71_294 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_71_283 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_44_497 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_176_108 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_158_812 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_157_300 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_161 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_150 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_194 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_183 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_172 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_8_321 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_145_517 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_138_591 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_141_712 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_125_274 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_113_425 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4270_ _7870_/Q _6486_/A1 _5849_/A2 _7572_/Q _4271_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_97_70 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_100_108 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_79_394 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_67_556 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_11_2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7960_ _7960_/D _7961_/RN _7960_/CLK _7960_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
X_7891_ _7891_/D _7901_/RN _7893_/CLK _7891_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
X_6911_ _6599_/Z _6941_/A2 _6908_/Z _7191_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor3_4
X_6842_ _7765_/Q _6892_/A2 _6892_/B1 _7731_/Q _6843_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_62_250 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_168_609 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_149_812 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3985_ _3985_/A1 _3985_/A2 _3985_/A3 _3985_/A4 _3990_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand4_1
X_6773_ _7656_/Q _6882_/B1 _6647_/Z _7616_/Q _6776_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_5724_ _5759_/A1 _5724_/A2 _5724_/B _5725_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_50_489 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_175_141 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_148_366 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_5655_ _5766_/A1 _5804_/A1 _5655_/A3 _5655_/A4 _5676_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor4_1
X_4606_ _4448_/Z _4608_/A2 _4606_/B _7405_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_7325_ _7901_/RN _4334_/Z _7325_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_117_753 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5586_ _5586_/A1 _5586_/A2 _5586_/A3 _5586_/A4 _5589_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand4_1
Xhold310 _7643_/Q hold310/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
X_4537_ _7377_/Q _4548_/A2 _4538_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
Xhold321 _7817_/Q hold321/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
XFILLER_116_263 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xhold343 _7691_/Q hold343/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
Xhold332 _7872_/Q hold332/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
X_7256_ _7256_/A1 _7256_/A2 _7257_/C VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_4468_ _7506_/Q _7263_/A1 hold40/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
Xhold387 _7797_/Q hold387/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
Xhold376 _7805_/Q hold376/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
Xhold354 _7707_/Q hold354/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
Xhold365 _7841_/Q hold365/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
X_6207_ hold349/Z _6208_/A2 _6208_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_104_469 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xhold398 _7370_/Q hold398/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
X_7187_ _7133_/S _7187_/A2 _7187_/B _7939_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_4399_ _7436_/Q input67/Z _7335_/Q _4399_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_86_810 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6138_ hold68/Z _6140_/A2 _6138_/B hold160/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_58_534 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_670 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_133_35 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_58_567 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_681 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_692 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_46_707 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6069_ hold393/Z _6072_/A2 _6070_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_18_409 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_26_33 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1825 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1814 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1803 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1858 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1847 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1836 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_81_570 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_54_795 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_158_108 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1869 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_41_467 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_53_294 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_179_480 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_182_612 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_158_87 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_154_325 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_139_388 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_5_302 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_182_667 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_181_144 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_135_561 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_123_712 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_5_357 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_174_64 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_107_296 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_150_575 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_123_778 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_122_266 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_95_128 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_67_73 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_49_567 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_64_526 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_49_578 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_29_280 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_44_250 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_177_428 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_60_743 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3770_ hold5/I _7968_/Q _3772_/S _7968_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_9_641 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5440_ _5705_/B _5712_/B _5555_/B _5534_/A2 _5444_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor4_1
XFILLER_8_195 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5371_ _5371_/A1 _5371_/A2 _5371_/B _5371_/C _5382_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_160_317 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_99_412 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_59_2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4322_ _4322_/A1 _4322_/A2 _7337_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_113_211 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7110_ _7714_/Q _7189_/A2 _7191_/B1 _7804_/Q _7111_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_113_233 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_7041_ _7833_/Q _7203_/A2 _6938_/I _7857_/Q _7043_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_4253_ _4253_/A1 _4253_/A2 _4253_/A3 _4253_/A4 _4263_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand4_1
XFILLER_101_428 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_99_489 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_86_117 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_86_128 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_95_651 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4184_ input47/Z _4231_/B1 _5817_/A1 _7559_/Q _5807_/A1 _7547_/Q _4186_/A1 VDD VSS
+ gf180mcu_fd_sc_mcu7t5v0__aoi222_1
Xclkbuf_3_4__f_wb_clk_i clkbuf_0_wb_clk_i/Z _7949_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_94_194 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_82_323 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7943_ _7943_/D _7949_/CLK _7943_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_55_537 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_82_389 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_63_570 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7874_ _7874_/D _7961_/RN _7874_/CLK _7874_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
X_6825_ _6825_/A1 _6825_/A2 _6825_/A3 _6826_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor3_1
X_3968_ _7827_/Q _6384_/A1 _3968_/B _3981_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_6756_ _7924_/Q _7133_/S _6757_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_5707_ _5782_/A2 _5704_/Z _5706_/Z _5717_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_164_601 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_149_686 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_148_174 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3899_ _7789_/Q _6299_/A1 _6435_/A1 _7853_/Q _3901_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_6687_ _7799_/Q _6883_/A2 _6883_/B1 _7783_/Q _6705_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_163_144 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_163_122 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5638_ _5064_/B _5678_/A3 _5637_/Z _7279_/B _5639_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai31_1
XFILLER_163_177 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5569_ _5376_/B _5218_/C _5587_/C VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_117_550 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_105_712 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xhold140 _7598_/Q hold140/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
Xhold162 hold162/I hold162/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
Xhold151 _7614_/Q hold151/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
X_7308_ input75/Z _4334_/Z _7308_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__and2_1
Xhold195 _7731_/Q hold195/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
Xhold173 hold173/I hold173/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
Xhold184 _7622_/Q hold184/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
X_7239_ _7518_/Q _7239_/A2 _7241_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_144_34 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_120_737 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_120_759 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_86_673 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_37_32 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_46_515 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2301 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_160_33 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2334 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2323 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2312 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1600 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2378 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2356 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2367 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2345 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_163_2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1633 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1622 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1611 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_61_529 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_26_250 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_2389 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1666 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1655 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1644 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_41_231 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_54_592 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_159_428 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1688 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1699 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1677 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_139_130 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_139_141 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_41_286 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_10_662 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_167_494 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_10_673 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_154_144 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_96_404 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_110_203 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_78_61 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_94_71 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_77_695 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_92_676 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_18_740 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4940_ _4946_/A1 _5230_/A1 _5200_/B _4974_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_4
XFILLER_64_389 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_45_570 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4871_ hold609/Z _4872_/A2 _4872_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_17_283 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_17_294 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3822_ _3801_/Z hold117/Z _3843_/A3 hold274/Z _4153_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand4_4
X_7590_ _7590_/D input75/Z _7889_/CLK _8000_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
X_6610_ _7434_/Q _7915_/Q _6610_/A3 _6611_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_177_269 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6541_ _4454_/Z _6553_/A2 _6541_/B _7895_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_146_601 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_145_100 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_3753_ _4383_/A1 _7413_/Q _4292_/B _3772_/S VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand3_4
XFILLER_173_442 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3684_ _7825_/Q _3684_/ZN VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_118_347 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6472_ hold639/Z _6485_/A2 _6473_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
Xoutput201 _4389_/ZN mgmt_gpio_oeb[37] VDD VSS gf180mcu_fd_sc_mcu7t5v0__buf_8
XFILLER_145_144 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5423_ _5624_/A1 _5648_/B2 _5724_/B _5627_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
Xoutput234 _4394_/Z mgmt_gpio_out[32] VDD VSS gf180mcu_fd_sc_mcu7t5v0__buf_8
XFILLER_145_177 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5354_ _5354_/A1 _5354_/A2 _5354_/A3 _5354_/A4 _5356_/A4 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor4_1
Xoutput212 _7989_/Z mgmt_gpio_out[12] VDD VSS gf180mcu_fd_sc_mcu7t5v0__buf_8
Xoutput223 _7996_/Z mgmt_gpio_out[22] VDD VSS gf180mcu_fd_sc_mcu7t5v0__buf_8
XFILLER_160_158 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4305_ _7414_/Q _4308_/S _7340_/Q _4306_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
Xoutput245 _4399_/Z mgmt_gpio_out[8] VDD VSS gf180mcu_fd_sc_mcu7t5v0__buf_8
Xoutput256 _4420_/ZN pad_flash_io1_oe VDD VSS gf180mcu_fd_sc_mcu7t5v0__buf_8
Xoutput267 _7556_/Q pll_ena VDD VSS gf180mcu_fd_sc_mcu7t5v0__buf_8
X_5285_ _5663_/A1 _5692_/B _5285_/A3 _5287_/C VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor3_1
XFILLER_101_203 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_99_286 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xoutput289 _7365_/Q pll_trim[2] VDD VSS gf180mcu_fd_sc_mcu7t5v0__buf_8
Xoutput278 _7347_/Q pll_trim[16] VDD VSS gf180mcu_fd_sc_mcu7t5v0__buf_8
X_7024_ _7816_/Q _7207_/A2 _7207_/B1 _7718_/Q _7024_/C _7025_/A4 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi221_1
X_4236_ _4236_/A1 _4236_/A2 _4236_/A3 _4236_/A4 _4283_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand4_2
XFILLER_114_37 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4167_ _4167_/A1 _4167_/A2 _4167_/A3 _4167_/A4 _4167_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__and4_1
X_4098_ _7750_/Q _6226_/A1 _6401_/A1 _7832_/Q _4100_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_7926_ _7926_/D _7961_/RN _7949_/CLK _7926_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_24_721 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7857_ _7857_/D _7901_/RN _7865_/CLK _7857_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
Xclkbuf_leaf_4_csclk clkbuf_leaf_9_csclk/I _7881_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
X_6808_ _7730_/Q _6892_/B1 _6880_/B1 _7812_/Q _6815_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_51_551 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_168_247 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7788_ _7788_/D _7901_/RN _7877_/CLK _7788_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_23_286 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_135_6 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6739_ _7647_/Q _6880_/C2 _6881_/B1 _7695_/Q _7809_/Q _6880_/B1 _6742_/A1 VDD VSS
+ gf180mcu_fd_sc_mcu7t5v0__aoi222_1
XFILLER_164_453 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_155_11 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_124_317 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_3_4 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_120_523 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_120_512 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_2_179 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_120_534 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_101_792 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_46_334 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_74_676 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_46_345 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_2153 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2142 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2131 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2120 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_27_570 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_46_389 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2186 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2175 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2164 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1441 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1430 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2197 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_159_203 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1474 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1452 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1463 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_120_91 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_120_80 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1496 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1485 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_14_275 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_128_656 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_127_133 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_127_144 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_6_463 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_123_361 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5070_ _5458_/C _5527_/A1 _5458_/B _5071_/C VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor3_1
XFILLER_111_556 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_97_779 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4021_ _7866_/Q _6469_/A1 _6418_/A1 _7842_/Q _4024_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_65_632 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5972_ hold643/Z _5987_/A2 _5973_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_80_602 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_64_175 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4923_ _4923_/A1 input97/Z _4926_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_7711_ _7711_/D _7901_/RN _7816_/CLK _7711_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_178_534 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_60_392 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4854_ hold659/Z _4857_/A2 _4855_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_7642_ _7642_/D _7961_/RN _7642_/CLK _7642_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_178_589 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_165_217 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3805_ hold116/Z _3803_/Z _3810_/S _3805_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_21_779 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7573_ _7573_/D input75/Z _7573_/CLK _7573_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
X_4785_ _7478_/Q _4795_/S _4786_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_3736_ _7976_/Q _3734_/Z _7978_/Q _3741_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_6524_ _4454_/Z _6536_/A2 _6524_/B _7887_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_118_166 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_3667_ hold14/I _7243_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_173_283 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6455_ hold640/Z _6468_/A2 _6456_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_5406_ _5292_/B _5779_/B1 _5587_/B _5406_/C _5407_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XFILLER_133_158 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6386_ _4448_/Z _6400_/A2 _6386_/B _7822_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_5337_ _5680_/A1 _5779_/A2 _5680_/B1 _5680_/B2 _5337_/C _5343_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi221_1
XFILLER_88_735 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_87_212 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_628 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_142_692 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5268_ _5394_/A1 _5005_/Z _5687_/B _5645_/A3 _5680_/C VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor4_2
XFILLER_141_180 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_125_47 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_102_534 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_87_223 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_125_69 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7007_ _7710_/Q _7189_/A2 _7191_/B1 _7800_/Q _7008_/A4 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_75_418 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_4219_ input11/Z _4219_/A2 _5812_/A1 _7556_/Q _4262_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_5199_ _4915_/Z _4996_/Z _5199_/B _5371_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_28_312 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_83_473 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_28_389 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_56_676 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_70_123 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_7909_ _7909_/D _7961_/RN _7940_/CLK _7909_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_4
XFILLER_24_573 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_34_33 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_169_567 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_157_707 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_11_212 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_8_717 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_126_2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_7_238 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_164_250 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_109_144 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_109_133 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_109_177 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_105_361 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_79_702 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_3_499 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_182_97 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_182_64 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_93_215 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_75_73 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_46_142 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_46_131 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_74_484 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_62_624 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_15_562 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1293 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1282 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1271 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1260 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_175_515 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_42_392 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4570_ hold720/Z _4573_/A2 _4571_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_156_751 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_155_283 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_116_615 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
Xhold728 _7741_/Q hold728/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
Xhold717 _7815_/Q hold717/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
XFILLER_7_783 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
Xhold706 hold706/I _5816_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
X_6240_ hold68/Z _6242_/A2 _6240_/B _7754_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_143_434 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_115_158 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_115_125 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
Xhold739 _7774_/Q hold739/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
X_6171_ hold277/Z _6174_/A2 _6172_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_41_2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5122_ _4953_/Z _5139_/A1 _5014_/Z _5122_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__and3_1
XFILLER_69_212 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_111_353 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_57_407 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5053_ _5199_/B _3727_/I _5303_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_4
X_4004_ _7890_/Q _6520_/A1 _4032_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_1_70 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_25_304 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_38_676 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_52_101 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_80_432 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_65_495 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5955_ hold743/Z _5970_/A2 _5956_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_4906_ _4905_/Z _5302_/A3 _4906_/S _4906_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_5886_ _5886_/A1 _7285_/A2 _5902_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_4
XFILLER_40_318 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_178_375 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4837_ _7519_/Q _7518_/Q _7520_/Q _5301_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__or3_1
X_7625_ _7625_/D _7961_/RN _7625_/CLK _7625_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
Xclkbuf_leaf_84_csclk _7558_/CLK _7876_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_146_250 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_7556_ _7556_/D input75/Z _7561_/CLK _7556_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
X_4768_ _4454_/Z _4768_/A2 _4768_/B hold580/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_4699_ _7988_/I _4718_/A1 _4702_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_106_103 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6507_ _4454_/Z _6519_/A2 _6507_/B _7879_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
Xclkbuf_leaf_99_csclk _7558_/CLK _7447_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
X_3719_ _7906_/Q _6633_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_3
X_7487_ _7487_/D _7912_/CLK _7487_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_162_743 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6438_ hold694/Z _6451_/A2 _6439_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_106_136 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_20_57 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_96_17 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_161_286 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_32
Xclkbuf_leaf_22_csclk _7825_/CLK _7809_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
X_6369_ _4448_/Z _6383_/A2 _6369_/B _7814_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_130_673 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_130_651 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xhold11 hold11/I hold11/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
Xhold22 hold22/I hold22/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
Xhold44 hold44/I hold44/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
Xhold55 hold55/I hold55/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
Xhold33 hold33/I hold33/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
XFILLER_75_215 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_29_77 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xhold88 hold88/I hold88/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
Xhold66 hold66/I hold66/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
Xhold99 hold99/I hold99/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
Xhold77 hold77/I hold77/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
Xclkbuf_leaf_37_csclk clkbuf_3_7__f_csclk/Z _7753_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_71_443 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_28_197 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_310 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_71_454 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_343 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_332 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_321 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
Xclkbuf_0_mgmt_gpio_in[4] mgmt_gpio_in[4] clkbuf_0_mgmt_gpio_in[4]/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_71_487 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XPHY_365 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_354 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_24_392 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_61_64 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_165_570 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_137_283 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_6_37 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_180_562 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_153_798 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_98_329 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_98_318 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_4_764 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_3_241 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_66_259 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_13_6 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_75_793 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_34_101 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_62_465 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_62_443 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_50_605 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_5740_ _5740_/A1 _5740_/A2 _5740_/A3 _5739_/Z _5804_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand4_1
XFILLER_15_381 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_22_318 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_22_329 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_148_504 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1090 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_5671_ _5774_/C _5671_/A2 _5748_/A2 _5671_/A4 _5671_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__or4_1
XFILLER_89_2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_7410_ _7410_/D _7901_/RN _7876_/CLK _7410_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
X_4622_ _3830_/Z _4448_/Z _4623_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_129_762 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_7341_ _7341_/D _7296_/Z _4031_/C2 _7341_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_128_250 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4553_ _4454_/Z _4553_/A2 _4553_/B _7384_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_7272_ _7272_/A1 _7280_/A2 _7277_/B _7272_/C _7273_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi211_1
X_4484_ _7506_/Q _7278_/A1 hold89/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_144_765 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xhold503 _7809_/Q hold503/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
Xhold525 _7899_/Q hold525/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
Xhold514 _7641_/Q hold514/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
Xhold536 hold536/I _4502_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
XFILLER_171_562 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6223_ hold68/Z _6225_/A2 _6223_/B _7746_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
Xhold547 hold547/I _7615_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
Xhold558 _7582_/Q hold558/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
Xhold569 _7404_/Q hold569/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
XFILLER_143_286 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_131_448 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6154_ hold280/Z _6157_/A2 _6155_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_830 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_841 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_852 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_6085_ hold47/Z _6089_/A2 _6085_/B _7681_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_112_673 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5105_ _5105_/A1 _5105_/A2 _5105_/A3 _5105_/A4 _5106_/A4 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand4_1
XTAP_863 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_874 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_885 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_57_215 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5036_ _5714_/A1 _5797_/A1 _5099_/B _5037_/C VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XTAP_896 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_122_37 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_26_602 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_25_167 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_41_605 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6987_ _7645_/Q _7195_/A2 _7195_/B1 _7621_/Q _7195_/C1 _7871_/Q _6990_/A2 VDD VSS
+ gf180mcu_fd_sc_mcu7t5v0__aoi222_1
X_5938_ hold767/Z _5953_/A2 _5939_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_40_126 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_179_673 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5869_ _7581_/Q hold26/Z hold27/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_7608_ _7608_/D _7961_/RN _7702_/CLK _7608_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_21_384 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_166_389 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7539_ _7539_/D _7959_/RN _7958_/CLK _7539_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_147_570 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_5_517 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_119_283 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_1_712 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xinput101 wb_adr_i[15] _4922_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_103_662 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_103_651 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_244 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_1_778 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
Xinput145 wb_dat_i[25] _7245_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
Xinput134 wb_dat_i[15] _7275_/B1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
Xinput112 wb_adr_i[25] _3660_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
Xinput123 wb_adr_i[6] _5199_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__buf_12
XFILLER_103_673 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_88_362 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
Xinput156 wb_dat_i[6] _7272_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_63_207 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_84_590 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_72_763 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_17_657 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_32_605 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_31_104 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_151 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_140 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
Xclkbuf_3_1__f_csclk clkbuf_0_csclk/Z clkbuf_leaf_9_csclk/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XPHY_184 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_173 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_162 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_9_812 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_145_507 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_195 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_172_326 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_172_348 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_180_392 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_140_212 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_125_286 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_99_638 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_141_779 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_140_256 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_79_340 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xclkbuf_3_3__f_wb_clk_i clkbuf_0_wb_clk_i/Z _7938_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_39_215 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_94_321 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_39_237 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_94_387 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_94_365 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7890_ _7890_/D _7901_/RN _7890_/CLK _7890_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_75_590 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6910_ _6599_/Z _6950_/A2 _6955_/A4 _7203_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor3_4
XFILLER_47_281 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6841_ _7829_/Q _6891_/A2 _6891_/B1 _7675_/Q _6891_/C1 _7781_/Q _6843_/A2 VDD VSS
+ gf180mcu_fd_sc_mcu7t5v0__aoi222_1
XFILLER_63_774 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_63_785 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_62_262 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_23_638 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3984_ _7713_/Q _6141_/A1 _6316_/A1 _7795_/Q _3985_/A4 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_6772_ _7648_/Q _6880_/C2 _6892_/A2 _7762_/Q _6776_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_5723_ _5723_/A1 _5723_/A2 _5791_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_176_676 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_5654_ _5740_/A3 _5651_/Z _5654_/A3 _5655_/A4 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_148_389 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_129_570 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4605_ hold715/Z _4608_/A2 _4606_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_7324_ _7901_/RN _4334_/Z _7324_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__and2_1
X_5585_ _5585_/A1 _5658_/B _5585_/B _5585_/C _5586_/A4 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi211_1
Xhold300 _8005_/I hold300/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
Xhold311 hold311/I _6004_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
X_4536_ _4454_/Z _4548_/A2 _4536_/B _7376_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
Xhold322 _7631_/Q hold322/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
Xhold333 _7719_/Q hold333/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
Xhold344 _7675_/Q hold344/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
X_7255_ _7520_/Q _7255_/A2 _7255_/B1 _7519_/Q _7256_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_1
Xhold377 _7690_/Q hold377/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
XFILLER_89_137 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xhold366 _7640_/Q hold366/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
X_4467_ _4487_/A1 hold73/Z _4467_/B hold482/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
Xhold355 _7578_/Q hold355/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
X_6206_ hold68/Z _6208_/A2 _6206_/B _7738_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_104_448 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4398_ _7437_/Q _4415_/A2 _7334_/Q _4398_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
Xhold388 _7802_/Q hold388/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
Xhold399 hold399/I _4521_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
X_7186_ _7939_/Q _7133_/S _7187_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_6137_ hold158/Z _6140_/A2 hold159/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_660 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_671 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_682 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_693 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_6068_ hold47/Z _6072_/A2 _6068_/B hold418/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_100_676 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_93_18 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_85_354 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5019_ _5200_/B _5230_/A1 _5024_/A2 _5201_/B _5021_/B1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai31_2
XFILLER_165_6 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1815 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1804 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_14_605 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_26_454 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1848 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1837 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1826 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_26_498 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_53_273 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1859 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_139_301 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_42_33 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_158_33 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_181_101 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_166_153 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_139_378 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_107_242 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_162_392 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_107_286 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_3_27 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_150_587 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_107_70 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_76_321 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_49_557 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_37_708 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_91_335 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_91_357 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_29_292 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_83_73 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_45_785 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_32_479 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_12_181 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_9_631 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_158_676 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_173_657 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_173_635 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5370_ _5369_/B _5381_/A2 _5370_/B _5375_/A4 VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_2
X_4321_ _4383_/A1 _7411_/Q _7337_/Q _4322_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_114_735 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_7040_ _7825_/Q _7202_/A2 _7201_/B1 _7671_/Q _7043_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_4252_ _7387_/Q _4559_/A1 _4779_/A1 _7476_/Q _4253_/A4 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_95_641 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4183_ _4183_/A1 _4183_/A2 _4183_/A3 _4187_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_94_151 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_67_354 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_27_207 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_103_39 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_7942_ _7942_/D _7944_/CLK _7942_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_36_730 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_36_741 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_7873_ _7873_/D _7901_/RN _7873_/CLK _7873_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_63_560 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_23_413 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_35_273 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_168_407 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6824_ _6824_/A1 _6824_/A2 _6824_/A3 _6824_/A4 _6825_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand4_1
XFILLER_63_593 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_23_424 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_35_295 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3967_ _4075_/B _4155_/A2 _3968_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_6755_ _7433_/Q _7923_/Q _6755_/B _6757_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_5706_ _5706_/A1 _5706_/A2 _5706_/A3 _5706_/A4 _5706_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__and4_1
XFILLER_50_298 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3898_ _7611_/Q _5920_/A1 _5971_/A1 _7635_/Q _3901_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_6686_ _7002_/B _6686_/A2 _6686_/A3 _6686_/B _7921_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai31_1
X_5637_ _5637_/A1 _5679_/A1 _5637_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_152_808 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5568_ _5104_/B _5708_/A2 _5578_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_151_318 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
Xhold130 _7342_/Q _3799_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
XFILLER_132_521 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xhold141 hold141/I _5909_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
XFILLER_88_29 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xhold152 hold152/I _7614_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
X_4519_ hold68/Z _4521_/A2 _4519_/B hold534/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_7307_ input75/Z _4334_/Z _7307_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__and2_1
X_7238_ _7279_/B _7238_/A2 _7238_/A3 _7280_/A3 _7277_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand4_4
X_5499_ _5499_/A1 _5499_/A2 _5653_/A1 _5499_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__or3_1
XFILLER_144_392 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xhold174 hold174/I _7440_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
Xhold163 hold163/I _7437_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
XFILLER_104_245 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
Xhold185 hold185/I _5960_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
XFILLER_144_57 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_104_278 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xhold196 _8000_/I hold196/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
XFILLER_58_321 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_7169_ _7535_/Q _7197_/A2 _7196_/A2 _7546_/Q _7196_/B1 _7474_/Q _7172_/A1 VDD VSS
+ gf180mcu_fd_sc_mcu7t5v0__aoi222_1
XTAP_490 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2302 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_100_484 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_100_495 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_100_473 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_46_549 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_2335 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2324 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2313 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_160_56 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_73_357 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_37_77 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_37_99 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2357 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2368 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2346 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1623 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1612 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1601 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_27_796 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2379 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_156_2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1667 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1656 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1645 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1634 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_744 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_53_32 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_1689 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1678 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_14_457 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_6_601 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_154_112 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_5_100 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_182_476 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_182_454 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_170_605 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_127_359 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_5_144 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_142_318 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_150_351 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_123_565 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_77_641 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_68_129 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_1_383 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_49_354 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_92_611 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_76_195 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_4870_ _4448_/Z _4872_/A2 _4870_/B _7527_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_32_210 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_177_226 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_177_215 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3821_ hold275/Z hold124/Z _6486_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_4
XFILLER_60_574 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6540_ hold589/Z _6553_/A2 _6541_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_33_799 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3752_ _3752_/I _3756_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_71_2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_146_646 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_118_337 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3683_ _7833_/Q _3683_/ZN VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_6471_ _4448_/Z _6485_/A2 _6471_/B _7862_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_9_494 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5422_ _5660_/A2 _5422_/A2 _5433_/C _5439_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
Xoutput235 _4395_/Z mgmt_gpio_out[33] VDD VSS gf180mcu_fd_sc_mcu7t5v0__buf_8
XFILLER_161_638 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_160_126 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xoutput213 _4412_/Z mgmt_gpio_out[13] VDD VSS gf180mcu_fd_sc_mcu7t5v0__buf_8
X_5353_ _5353_/A1 _5642_/A2 _5493_/B _5353_/A4 _5354_/A4 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand4_1
Xoutput224 _7997_/Z mgmt_gpio_out[23] VDD VSS gf180mcu_fd_sc_mcu7t5v0__buf_8
XFILLER_99_210 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
Xoutput202 _3709_/ZN mgmt_gpio_oeb[3] VDD VSS gf180mcu_fd_sc_mcu7t5v0__buf_8
X_4304_ _4304_/I0 _7342_/Q _4309_/S _7342_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_126_392 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xoutput246 _4398_/Z mgmt_gpio_out[9] VDD VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
Xoutput268 _7563_/Q pll_sel[0] VDD VSS gf180mcu_fd_sc_mcu7t5v0__buf_8
Xoutput257 _7566_/Q pll90_sel[0] VDD VSS gf180mcu_fd_sc_mcu7t5v0__buf_8
XFILLER_141_351 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5284_ _5573_/A1 _5292_/B _5247_/B _5431_/B _5288_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_1
Xoutput279 _7348_/Q pll_trim[17] VDD VSS gf180mcu_fd_sc_mcu7t5v0__buf_8
X_7023_ _7023_/A1 _7023_/A2 _7023_/A3 _7024_/C VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_101_215 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_4235_ _7822_/Q _6384_/A1 _4863_/A1 _7525_/Q _4236_/A4 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_4166_ _7364_/Q _4505_/A1 _6005_/A1 _7645_/Q _4167_/A4 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_28_527 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4097_ _7654_/Q _6022_/A1 _6537_/A1 _7896_/Q _4100_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_55_357 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_82_176 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7925_ _7925_/D _7961_/RN _7938_/CLK _7925_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_169_716 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_130_37 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_7856_ _7856_/D _7901_/RN _7890_/CLK _7856_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffsnq_1
XFILLER_23_210 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_24_744 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6807_ _7796_/Q _6893_/A2 _6890_/B1 _7852_/Q _6815_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_168_259 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4999_ _4999_/A1 _4999_/A2 _4999_/A3 _4999_/A4 _4999_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__and4_1
X_7787_ _7787_/D _7901_/RN _7901_/CLK _7787_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
X_6738_ _6738_/A1 _6738_/A2 _6738_/A3 _6738_/A4 _6753_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand4_1
XFILLER_109_337 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6669_ _7822_/Q _6891_/A2 _6894_/C1 _7830_/Q _6683_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_152_605 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_155_23 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_136_189 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_117_381 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_105_532 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_59_641 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_93_408 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_86_460 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_86_471 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_58_173 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2110 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_104_60 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_73_121 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2143 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2132 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2121 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_34_519 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2176 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2165 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2154 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1442 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1431 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1420 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_73_198 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_2198 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2187 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_159_215 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1475 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1453 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1464 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_14_254 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_159_237 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1497 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1486 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_15_799 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_30_747 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_128_602 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_155_421 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_128_646 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_10_460 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_127_156 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_155_487 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_143_638 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_142_104 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_115_318 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_108_392 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_151_682 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_97_747 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_111_579 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_84_419 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4020_ _4020_/A1 _4020_/A2 _4020_/A3 _4020_/A4 _4025_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand4_1
XFILLER_49_140 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_49_173 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_92_441 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_64_143 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_64_132 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_37_357 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5971_ _5971_/A1 hold32/Z _5987_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_4
XFILLER_92_463 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_25_519 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4922_ input99/Z input98/Z _4922_/A3 _4922_/A4 _4926_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand4_1
X_7710_ _7710_/D _7901_/RN _7753_/CLK _7710_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffsnq_1
X_7641_ _7641_/D _7961_/RN _7649_/CLK _7641_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
X_4853_ _4853_/A1 _7285_/A2 _4857_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_3804_ _7506_/Q hold116/Z _3806_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__and2_1
X_4784_ _7515_/Q _7959_/RN _4795_/S VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_4
XFILLER_21_758 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7572_ _7572_/D _7572_/CLK _7572_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffq_1
Xclkbuf_opt_2_0_csclk clkbuf_3_6__f_csclk/Z clkbuf_opt_2_0_csclk/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
X_3735_ _4380_/B _3734_/Z _3735_/B _7979_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_6523_ hold594/Z _6536_/A2 _6524_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_174_763 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_134_605 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_109_16 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6454_ _4448_/Z _6468_/A2 _6454_/B _7854_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_5405_ _5701_/A2 _5682_/A3 _5405_/B _5406_/C VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_106_318 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_133_137 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_127_690 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_6385_ hold742/Z _6400_/A2 _6386_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_5336_ _5394_/A1 _5344_/A2 _5687_/B _5618_/A3 _5337_/C VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor4_1
X_5267_ _5433_/C _5573_/A1 _5722_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_88_747 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7006_ _7686_/Q _7189_/B1 _7189_/C1 _7654_/Q _7008_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_4218_ _7782_/Q _6299_/A1 _6248_/A1 _7758_/Q _4262_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_5198_ _5015_/B _5371_/C _5197_/Z _7519_/Q _5415_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai31_2
XFILLER_68_471 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_44_806 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4149_ _4153_/A1 _3881_/Z _4774_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_55_121 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_28_379 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_83_496 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_24_530 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7908_ _7908_/D _7961_/RN _7940_/CLK _7908_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_4
XFILLER_70_168 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_70_157 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_70_179 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_7839_ _7839_/D input75/Z _7886_/CLK _7839_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffsnq_1
XFILLER_12_747 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_24_596 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_149_270 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_50_33 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_166_33 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_109_156 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_165_785 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_152_402 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_125_638 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_124_104 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_119_2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_180_744 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_118_690 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_152_479 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_124_159 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_1_2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_120_321 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_105_384 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_182_76 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_87_791 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_87_780 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_59_482 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_74_441 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_19_357 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_74_463 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_46_176 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1250 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_91_73 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_1283 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1272 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1261 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_70_680 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1294 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_116_605 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_11_780 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_115_104 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
Xhold707 hold707/I _7557_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
XFILLER_6_250 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xhold718 _7653_/Q hold718/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
Xhold729 _7791_/Q hold729/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
XFILLER_131_619 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_6170_ hold47/Z _6174_/A2 _6170_/B _7721_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_5121_ _5087_/B _5680_/B2 _5218_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
Xclkbuf_leaf_3_csclk clkbuf_leaf_9_csclk/I _7890_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_34_2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5052_ _5452_/C _5543_/C _5797_/A2 _5064_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor3_2
XFILLER_111_365 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_84_238 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4003_ _7874_/Q _6486_/A1 _4035_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_37_110 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_93_783 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_1_82 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5954_ _5954_/A1 _7285_/A2 _5970_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_4
XFILLER_178_332 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_178_321 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4905_ _5224_/A3 _5224_/A4 _4905_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__and2_1
X_5885_ _4454_/Z _5885_/A2 _5885_/B _7587_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_52_179 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4836_ _7519_/Q _7518_/Q _7520_/Q _7280_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor3_4
X_7624_ _7624_/D _7961_/RN _7642_/CLK _7624_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
X_7555_ _7555_/D _7314_/Z _4418_/I1 _7555_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffnrnq_1
XFILLER_147_763 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6506_ hold655/Z _6519_/A2 _6507_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_4767_ hold579/Z _4768_/A2 _4768_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_4698_ _4718_/A1 _4698_/A2 _4698_/B hold171/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_112_9 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_107_638 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3718_ _7907_/Q _6634_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__inv_2
X_7486_ _7486_/D _7912_/CLK _7486_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_6437_ _4448_/Z _6451_/A2 _6437_/B _7846_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_3649_ _7903_/Q _6565_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_6368_ hold766/Z _6383_/A2 _6369_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_136_69 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5319_ _5563_/B2 _5365_/B1 _5319_/B _5319_/C _5419_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi211_4
XFILLER_121_129 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_121_118 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_114_170 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_102_321 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xhold23 hold23/I hold23/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
Xhold12 hold12/I hold12/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
X_6299_ _6299_/A1 _7285_/A2 _6315_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_4
Xhold45 hold45/I hold45/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
Xhold34 hold34/I hold34/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
Xhold56 hold56/I hold56/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
XFILLER_130_696 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_69_780 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xhold67 hold67/I hold67/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
Xhold89 hold89/I hold89/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
Xhold78 hold78/I hold78/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
XFILLER_91_709 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_28_132 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_16_305 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_56_463 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_71_422 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_28_176 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_300 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_45_66 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_169_343 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_333 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_322 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_311 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_71_499 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XPHY_355 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_177_10 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_344 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_169_354 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_61_98 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_152_276 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_3_231 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_106_671 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_3_286 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_121_641 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xclkbuf_3_2__f_wb_clk_i clkbuf_0_wb_clk_i/Z _7940_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_67_728 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_75_783 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_62_433 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_62_411 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_34_157 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_34_179 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_5670_ _5799_/A1 _5799_/A2 _5776_/A4 _5799_/A3 _5671_/A4 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand4_1
XTAP_1091 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1080 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_4621_ _7990_/I _4652_/A1 _4624_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_175_357 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_7340_ _7340_/D _7295_/Z _4415_/A2 _7340_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_129_785 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_116_402 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4552_ hold612/Z _4553_/A2 _4553_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_7271_ _7271_/A1 _7271_/A2 _7272_/C VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_144_744 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xhold504 _7900_/Q hold504/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
Xhold526 _8003_/I hold526/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
Xhold515 hold515/I _7641_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
XFILLER_7_570 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4483_ hold297/Z _4487_/A1 hold298/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_6222_ hold437/Z _6225_/A2 _6223_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
Xhold559 _7457_/Q hold559/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
Xhold548 _7366_/Q hold548/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
Xhold537 hold537/I _7361_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
XFILLER_131_416 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_103_129 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_103_118 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6153_ hold47/Z _6157_/A2 _6153_/B _7713_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
XTAP_820 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_831 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_842 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_853 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_6084_ hold412/Z _6089_/A2 _6085_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_112_685 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5104_ _5705_/A2 _5783_/A2 _5104_/B _5105_/A4 VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_85_503 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_864 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_875 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_886 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_5035_ _5069_/A2 _4930_/Z _4953_/Z _5035_/A4 _5099_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand4_4
XFILLER_111_184 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_73_709 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_897 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_38_463 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_25_102 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6986_ _6986_/A1 _6986_/A2 _6991_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_179_641 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_81_797 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5937_ _5937_/A1 hold32/Z _5953_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_4
XFILLER_40_105 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_53_499 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_178_151 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5868_ _4454_/Z _5868_/A2 _5868_/B _7580_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_7607_ _7607_/D _7961_/RN _7645_/CLK _7607_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffsnq_2
XFILLER_21_363 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_5799_ _5799_/A1 _5799_/A2 _5799_/A3 _5799_/A4 _5800_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand4_1
X_4819_ _7219_/A1 _4828_/S _4819_/B _7496_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_7538_ _7538_/D _7961_/RN _7960_/CLK _7538_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_134_232 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7469_ _7469_/D _7961_/RN _7532_/CLK _7469_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_135_766 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_150_747 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_212 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xinput102 wb_adr_i[16] _4924_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_163_23 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_103_641 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_1_757 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_49_706 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xinput135 wb_dat_i[16] _7239_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
Xinput124 wb_adr_i[7] _3727_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_12
Xinput113 wb_adr_i[26] _3661_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_130_460 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_76_514 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
Xinput146 wb_dat_i[26] _7250_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
Xinput157 wb_dat_i[7] _7277_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_76_547 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_91_539 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_84_580 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_29_496 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_44_411 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_44_422 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_57_783 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_16_179 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_44_477 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_169_140 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_152 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_141 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_130 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_157_313 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_185 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_174 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_163 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_157_357 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_196 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_165_390 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_126_744 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_98_105 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_95_812 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xclkbuf_leaf_83_csclk clkbuf_leaf_9_csclk/I _7582_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_67_547 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_63_720 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6840_ _7797_/Q _6893_/A2 _6893_/B1 _7773_/Q _6893_/C1 _7635_/Q _6843_/A1 VDD VSS
+ gf180mcu_fd_sc_mcu7t5v0__aoi222_1
XFILLER_90_550 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_63_764 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_62_241 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6771_ _6771_/A1 _6771_/A2 _6771_/A3 _6771_/A4 _6777_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand4_1
XFILLER_22_105 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_23_628 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_35_499 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5722_ _5722_/A1 _5620_/B _5722_/B _5723_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_3983_ _7352_/Q _4444_/A1 _4505_/A1 _7368_/Q _3985_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_1
Xclkbuf_leaf_21_csclk _7825_/CLK _7851_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
X_5653_ _5653_/A1 _5542_/Z _5764_/A2 _5746_/A4 _5654_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor4_1
X_5584_ _5704_/A1 _5716_/A2 _5732_/A2 _5794_/A2 _5589_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand4_1
X_4604_ _4604_/A1 _7285_/A2 _4608_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
Xhold301 _7378_/Q hold301/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
X_4535_ hold690/Z _4548_/A2 _4536_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
Xclkbuf_leaf_36_csclk clkbuf_3_7__f_csclk/Z _7813_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
X_7323_ _7901_/RN _4334_/Z _7323_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_7_70 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xhold334 _7850_/Q hold334/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
Xhold323 hold323/I _7631_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
XFILLER_117_16 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
Xhold312 hold312/I _7643_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
X_7254_ _7518_/Q _7254_/A2 _7256_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_132_747 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_132_725 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
Xhold345 hold345/I _7675_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
Xhold378 _7610_/Q hold378/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
Xhold367 hold367/I _7640_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
X_4466_ hold480/Z _4487_/A1 hold481/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
Xhold356 _7624_/Q hold356/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
Xhold389 _7738_/Q hold389/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
X_6205_ hold389/Z _6208_/A2 _6206_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_4397_ _7438_/Q input58/Z _7335_/Q _4397_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_7185_ _7433_/Q _7938_/Q _7185_/B _7187_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_112_460 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_112_471 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6136_ hold47/Z _6140_/A2 _6136_/B _7705_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_97_160 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_86_812 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_58_525 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_650 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_661 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_58_558 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_672 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_683 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_694 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_6067_ hold417/Z _6072_/A2 _6068_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_46_709 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5018_ _5529_/A2 _5529_/A3 _5528_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_2
XFILLER_26_411 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_39_783 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_39_794 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1816 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1805 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1849 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1838 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1827 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_14_617 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_41_414 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_53_252 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_6969_ _7846_/Q _7193_/A2 _7205_/A2 _7732_/Q _6971_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_41_425 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_179_482 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_167_611 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_10_801 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_139_357 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_21_171 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_166_176 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_127_519 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_108_744 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_108_788 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_101_2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_174_33 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_122_213 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_77_812 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_1_565 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_49_514 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_131_780 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_49_525 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_76_388 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_72_550 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_45_742 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_17_499 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_32_447 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_32_458 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_32_469 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_157_110 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_9_621 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_157_187 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_172_179 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4320_ _7336_/Q _4300_/C _4322_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_126_585 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_99_425 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_114_747 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_99_447 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_4_392 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4251_ _7644_/Q _6005_/A1 _4883_/A1 _7533_/Q _4253_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_101_408 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_86_108 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_86_119 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_68_812 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4182_ _7693_/Q _6107_/A1 _4858_/A1 _7524_/Q _4183_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_7941_ _7941_/D _7959_/RN _7958_/CLK _7941_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_103_29 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_7872_ _7872_/D _7901_/RN _7899_/CLK _7872_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffsnq_1
XFILLER_51_712 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6823_ _7714_/Q _6885_/B1 _6890_/A2 _7642_/Q _6824_/A4 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_23_436 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_50_211 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3966_ _7673_/Q _6056_/A1 _5937_/A1 _7617_/Q _3992_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_6754_ _6754_/A1 _6767_/C _6754_/B1 _6754_/B2 _7433_/Q _6755_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi221_1
XFILLER_51_778 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5705_ _5104_/B _5705_/A2 _5705_/B _5706_/A4 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_10_108 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_6685_ _7604_/Q _7910_/Q _6879_/A1 _6686_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor3_1
XFILLER_176_463 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5636_ _5636_/A1 _5417_/I _5708_/B _5679_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor3_1
X_3897_ _7755_/Q _6226_/A1 _6401_/A1 _7837_/Q _3901_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_163_113 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_148_176 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_128_37 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_12_37 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_128_48 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_117_552 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5567_ _4998_/B _5412_/B _5567_/A3 _5706_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor3_1
Xhold120 hold120/I _7726_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
X_5498_ _5689_/A2 _5498_/A2 _5498_/B _5543_/C _5653_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi211_1
Xhold131 hold131/I hold131/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
Xhold153 _7336_/Q hold153/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
Xhold142 hold142/I _7598_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
X_4518_ hold532/Z _4521_/A2 hold533/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_2_318 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7306_ input75/Z _4334_/Z _7306_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__and2_1
X_7237_ _7516_/Q _7237_/A2 _7280_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_4449_ hold15/Z _4449_/A2 hold16/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
Xhold164 _7596_/Q hold164/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
XFILLER_105_769 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
Xhold175 _7638_/Q hold175/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
Xhold186 hold186/I _7622_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
Xhold197 _7996_/I hold197/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
XFILLER_120_717 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_59_812 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_132_599 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_113_780 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7168_ _7168_/A1 _7168_/A2 _7178_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_7099_ _7737_/Q _7205_/A2 _7205_/B1 _7745_/Q _7100_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_6119_ hold47/Z _6123_/A2 _6119_/B _7697_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
XTAP_491 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_480 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_19_709 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_100_463 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_58_388 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2325 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2314 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2303 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_160_68 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2369 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2347 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2358 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2336 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_163_4 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_160_79 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1624 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1613 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1602 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1657 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1646 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1635 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_14_447 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_149_2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1679 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1668 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_767 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_167_430 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_139_132 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_22_480 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_139_154 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_182_422 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_167_496 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_127_327 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_10_664 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_154_157 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_182_499 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_182_488 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_154_179 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_5_167 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_5_156 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_150_330 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xclkbuf_1_0__f__1040_ clkbuf_0__1040_/Z _4807_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_111_728 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_111_706 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_68_108 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_68_119 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_1_373 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_76_141 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_91_144 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_64_358 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_92_689 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_33_712 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_91_188 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_3820_ hold123/Z _3925_/A2 _3790_/Z _3963_/A4 hold124/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand4_4
XFILLER_60_586 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_20_439 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_32_299 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3751_ _3730_/Z _3751_/A2 _3751_/A3 _3752_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor3_1
XFILLER_158_463 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3682_ _7841_/Q _3682_/ZN VDD VSS gf180mcu_fd_sc_mcu7t5v0__inv_1
X_6470_ hold732/Z _6485_/A2 _6471_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_9_473 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5421_ _5421_/A1 _5421_/A2 _5421_/A3 _5421_/B1 _5498_/A2 _5422_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai32_1
XFILLER_133_308 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_64_2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_173_499 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_160_105 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xoutput214 _4411_/Z mgmt_gpio_out[14] VDD VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
Xoutput225 _7998_/Z mgmt_gpio_out[24] VDD VSS gf180mcu_fd_sc_mcu7t5v0__buf_8
X_5352_ _5788_/A2 _5534_/A2 _5353_/A4 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_1
Xoutput203 _3708_/ZN mgmt_gpio_oeb[4] VDD VSS gf180mcu_fd_sc_mcu7t5v0__buf_8
Xoutput236 _8006_/Z mgmt_gpio_out[34] VDD VSS gf180mcu_fd_sc_mcu7t5v0__buf_8
X_4303_ _7414_/Q _4297_/Z _4303_/A3 _4303_/B _4304_/I0 VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai31_1
XFILLER_141_330 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_114_544 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
Xoutput258 _7567_/Q pll90_sel[1] VDD VSS gf180mcu_fd_sc_mcu7t5v0__buf_8
Xoutput247 _4418_/Z pad_flash_clk VDD VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
X_7022_ _7734_/Q _7205_/A2 _7205_/B1 _7742_/Q _7023_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_5283_ _5247_/B _5624_/B _5783_/B _5288_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_87_417 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_87_428 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xoutput269 _7564_/Q pll_sel[1] VDD VSS gf180mcu_fd_sc_mcu7t5v0__buf_8
X_4234_ _7604_/Q _5920_/A1 _4873_/A1 _7529_/Q _4236_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_68_664 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_67_141 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_67_130 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4165_ _7815_/Q hold134/I _4609_/A1 _7408_/Q _4843_/A1 _7508_/Q _4167_/A3 VDD VSS
+ gf180mcu_fd_sc_mcu7t5v0__aoi222_1
XFILLER_95_494 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_83_623 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_67_152 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4096_ _7377_/Q hold114/I _4239_/A2 input22/Z hold108/I input63/Z _4100_/A1 VDD VSS
+ gf180mcu_fd_sc_mcu7t5v0__aoi222_1
X_7924_ _7924_/D _7961_/RN _7938_/CLK _7924_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
X_7855_ _7855_/D _7901_/RN _7890_/CLK _7855_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffsnq_1
XFILLER_36_594 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6806_ _7706_/Q _6889_/A2 _6805_/Z _6830_/B _6819_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_24_789 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4998_ _5705_/A2 _4996_/Z _4998_/B _4998_/C _4999_/A4 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi211_1
X_7786_ _7786_/D _7901_/RN _7881_/CLK _7786_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_11_428 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_177_783 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_164_400 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_135_8 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6737_ _7793_/Q _6893_/A2 _6893_/B1 _7769_/Q _6738_/A4 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_3949_ input59/Z _5886_/A1 _4219_/A2 input18/Z _6469_/A1 _7868_/Q _3953_/A1 VDD VSS
+ gf180mcu_fd_sc_mcu7t5v0__aoi222_2
XFILLER_176_282 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_149_485 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_139_69 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6668_ _7375_/Q _6882_/A2 _6665_/Z _7740_/Q _6683_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_136_135 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5619_ _5319_/C _5714_/B1 _5319_/B _5619_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__or3_1
X_6599_ _7912_/Q _6599_/A2 _6599_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__or2_4
XFILLER_136_179 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_155_57 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_3_638 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_48_33 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_120_569 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_101_783 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_100_271 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_46_314 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2100 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_73_144 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_58_185 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2144 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2133 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2111 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2122 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_64_54 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_15_712 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2177 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2166 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2155 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1432 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1421 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1410 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_531 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2199 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2188 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_159_205 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1454 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1465 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1443 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_542 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_175_709 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1498 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1487 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1476 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_14_277 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_30_759 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_127_113 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_127_124 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_80_97 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_155_444 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_182_274 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_155_499 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_142_116 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_127_168 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_89_73 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_69_428 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_96_247 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_77_494 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_37_347 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_53_807 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5970_ hold90/Z _5970_/A2 _5970_/B hold309/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_25_509 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4921_ _4917_/Z _4919_/Z _5210_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_4
XFILLER_80_637 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4852_ _4454_/Z _4852_/A2 _4852_/B hold603/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_7640_ _7640_/D _7961_/RN _7643_/CLK _7640_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_33_553 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_33_564 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3803_ hold753/Z hold628/Z _7414_/Q _3803_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_4783_ _4454_/Z _4783_/A2 _4783_/B hold598/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_7571_ _7571_/D _7961_/RN _7625_/CLK _7571_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffsnq_1
XFILLER_159_783 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_158_282 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_146_422 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_118_102 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6522_ _4448_/Z _6536_/A2 _6522_/B _7886_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_3734_ _7414_/Q _7413_/Q _7411_/Q _3734_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__or3_2
XFILLER_109_28 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3665_ _7607_/Q _6754_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_6453_ hold731/Z _6468_/A2 _6454_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_161_425 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5404_ _5404_/A1 _5779_/B1 _5682_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_133_105 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_118_179 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6384_ _6384_/A1 _7285_/A2 _6400_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_4
XFILLER_142_672 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5335_ _5335_/A1 _5335_/A2 _5331_/Z _5335_/A4 _5354_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand4_1
XFILLER_130_812 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_142_694 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5266_ _5687_/B _5645_/A3 _5680_/B1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_141_193 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7005_ _7678_/Q _7191_/A2 _7190_/B1 _7614_/Q _7190_/A2 _7792_/Q _7008_/A2 VDD VSS
+ gf180mcu_fd_sc_mcu7t5v0__aoi222_1
X_4217_ hold275/Z _4217_/A2 _5871_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_5197_ _5209_/A2 _5209_/A3 _5197_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__and2_1
X_4148_ _4153_/A1 hold156/Z _4764_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_55_133 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_4079_ _7662_/Q _6039_/A1 _6452_/A1 _7856_/Q _4080_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_55_144 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_71_659 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_71_637 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_70_103 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7907_ _7907_/D _7961_/RN _7940_/CLK _7907_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffsnq_4
XFILLER_169_503 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7838_ _7838_/D _7901_/RN _7881_/CLK _7838_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffsnq_1
XFILLER_12_737 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_157_709 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7769_ _7769_/D _7901_/RN _7890_/CLK _7769_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_137_422 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_164_263 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_137_499 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_109_179 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_109_168 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_180_767 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_117_190 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_105_341 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_182_33 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_78_203 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_59_65 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xclkbuf_3_1__f_wb_clk_i clkbuf_0_wb_clk_i/Z _7944_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_78_258 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_78_247 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_59_450 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_101_580 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_59_494 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_19_369 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_34_306 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_46_166 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_62_637 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1240 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1284 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1273 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1262 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1251 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_15_586 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1295 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_30_534 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_30_523 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_42_383 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_147_219 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_11_770 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_128_433 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_171_712 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
Xhold708 _7871_/Q hold708/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
Xhold719 _7385_/Q hold719/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
XFILLER_170_211 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_143_425 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_115_116 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_6_273 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_130_108 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_124_661 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_112_812 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5120_ _5319_/C _5689_/A2 _5390_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_123_160 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_97_523 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_97_512 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5051_ _5006_/C _5448_/A1 _5797_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_4
XFILLER_123_182 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_97_567 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_27_2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_97_589 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4002_ _4002_/A1 _4427_/B _4002_/B1 _4002_/B2 _7553_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_92_250 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_65_475 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_37_144 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_53_626 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_53_648 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_179_812 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5953_ hold90/Z _5953_/A2 _5953_/B hold352/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_80_456 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4904_ _5087_/C _4900_/Z _5496_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_4
X_5884_ hold619/Z _5885_/A2 _5885_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_33_350 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_166_517 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_139_709 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7623_ _7623_/D _7961_/RN _7649_/CLK _7623_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
X_4835_ _4454_/Z _4835_/A2 _4835_/B hold623/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_147_720 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4766_ _4448_/Z _4768_/A2 _4766_/B _7470_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_21_567 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7554_ _7554_/D _7313_/Z _7977_/CLK _7554_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffnrnq_1
X_6505_ _4448_/Z _6519_/A2 _6505_/B _7878_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_3717_ _7910_/Q _6878_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_12
XFILLER_162_723 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_134_414 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4697_ hold140/Z _3819_/Z _4697_/B _4698_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_106_105 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7485_ _7485_/D _7944_/CLK _7485_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_6436_ hold760/Z _6451_/A2 _6437_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_119_499 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_106_138 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_20_37 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3648_ _7432_/Q _6572_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_136_37 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6367_ hold134/Z hold32/Z _6383_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_4
X_5318_ _5350_/A3 _5495_/B2 _5555_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_2
XFILLER_103_812 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_88_534 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6298_ hold90/Z _6298_/A2 _6298_/B _7781_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_88_545 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
Xhold13 hold13/I hold13/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
XFILLER_0_449 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xhold35 hold35/I hold35/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
Xhold46 hold46/I hold46/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
X_5249_ _3728_/I _5022_/B _5054_/Z _5687_/B _5425_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor4_4
Xhold24 hold24/I hold24/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
Xhold79 hold79/I hold79/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
Xhold68 hold68/I hold68/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
Xhold57 hold57/I hold57/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
XFILLER_28_122 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_29_634 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_56_453 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_83_283 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_301 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_71_456 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_334 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_323 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_312 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_40_810 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_356 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_345 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_101_73 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_12_534 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_12_523 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_169_377 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_131_2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_129_219 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_8_527 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_153_712 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_180_531 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_152_200 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_152_211 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_125_425 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_4_733 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_180_564 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_152_255 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_140_417 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_112_119 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_112_108 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_79_567 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_67_707 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_120_152 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_39_409 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_81_209 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_74_250 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_19_144 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_90_743 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_34_169 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_1092 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1081 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1070 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_175_303 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4620_ _4620_/A1 _5903_/A2 _4686_/B1 _3830_/Z hold12/Z _4652_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi221_4
XFILLER_129_720 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4551_ _4448_/Z _4553_/A2 _4551_/B _7383_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_7270_ _7520_/Q _7270_/A2 _7270_/B1 _7518_/Q _7271_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_1
Xhold505 _7884_/Q hold505/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
Xhold516 _7859_/Q hold516/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
X_4482_ _4487_/A1 hold68/Z _4482_/B hold432/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
Xhold527 _7623_/Q hold527/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
X_6221_ hold47/Z _6225_/A2 _6221_/B hold271/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_143_244 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_131_406 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
Xhold538 _7833_/Q hold538/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
Xhold549 hold549/I _4513_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
X_6152_ hold284/Z _6157_/A2 _6153_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_131_428 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_810 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_5103_ _5669_/B _5669_/A1 _5648_/A2 _5104_/B _5105_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XTAP_821 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_832 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_843 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_111_141 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_100_804 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_97_375 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6083_ hold41/Z _6089_/A2 _6083_/B _7680_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
XTAP_854 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_865 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_876 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_5034_ _5661_/A1 _4965_/B _5647_/A2 _5752_/B1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor3_4
XTAP_887 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_898 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_38_453 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_93_570 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_65_283 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_65_294 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6985_ _7693_/Q _7194_/A2 _7194_/B1 _7661_/Q _7194_/C1 _7807_/Q _6986_/A2 VDD VSS
+ gf180mcu_fd_sc_mcu7t5v0__aoi222_1
XFILLER_53_456 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5936_ hold90/Z _5936_/A2 _5936_/B _7611_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_22_810 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_25_169 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_178_174 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7606_ _7606_/D _7961_/RN _7702_/CLK _7606_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
X_5867_ hold564/Z _5868_/A2 _5868_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_182_807 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_166_347 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_119_230 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5798_ _5583_/C _5185_/B _5798_/A3 _5798_/A4 _5799_/A4 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor4_1
X_4818_ _7496_/Q _4828_/S _4819_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_4749_ hold641/Z _4749_/I1 _4753_/S _7462_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_147_561 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_135_712 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_119_241 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_7537_ _7537_/D _7961_/RN _7642_/CLK _7537_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_134_211 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_107_425 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7468_ _7468_/D _7961_/RN _7532_/CLK _7468_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
X_6419_ hold733/Z _6434_/A2 _6420_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_7399_ _7399_/D _7961_/RN _7756_/CLK _7399_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_1_769 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
Xinput136 wb_dat_i[17] _7244_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
Xinput114 wb_adr_i[27] _4368_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
Xinput103 wb_adr_i[17] _4924_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
Xinput125 wb_adr_i[8] _4923_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_102_152 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_279 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_49_729 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xinput147 wb_dat_i[27] _7255_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
Xinput158 wb_dat_i[8] _7240_/B1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_102_174 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_29_442 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_56_33 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_179_2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_56_250 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_112_50 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_71_231 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_16_136 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_112_83 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_112_72 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_44_489 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_71_286 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XPHY_142 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_131 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_120 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_31_117 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_175 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
Xclkbuf_leaf_2_csclk clkbuf_leaf_9_csclk/I _7865_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XPHY_164 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_153 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_24_191 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_169_196 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_197 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_186 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_40_673 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_125_211 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_125_233 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_113_417 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_113_428 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_98_128 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_140_247 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_98_139 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_97_73 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_97_62 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_94_301 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_67_515 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_48_740 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_94_389 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_82_529 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_75_592 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_75_570 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_35_423 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_47_283 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3982_ _7851_/Q _6435_/A1 _6469_/A1 _7867_/Q _3985_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_90_562 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6770_ _7818_/Q _6880_/A2 _6893_/C1 _7632_/Q _6771_/A4 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XPHY_0 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_149_804 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5721_ _5621_/B _5724_/A2 _5721_/B _5721_/C _5722_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XFILLER_94_2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_175_100 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_50_459 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5652_ _5162_/B _5652_/A2 _5652_/A3 _5652_/A4 _5746_/A4 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand4_1
XFILLER_148_325 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_175_155 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_175_144 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_129_561 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_117_712 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5583_ _5062_/Z _5690_/A1 _5583_/B _5583_/C _5794_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi211_1
X_4603_ _4454_/Z _4603_/A2 _4603_/B _7404_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_7322_ _7901_/RN _4334_/Z _7322_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__and2_1
Xhold302 _7752_/Q hold302/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
XFILLER_156_380 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_4534_ _4448_/Z _4548_/A2 _4534_/B _7375_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_144_531 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_116_200 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
Xhold324 _7832_/Q hold324/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
Xhold335 _8004_/I hold335/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
X_7253_ _7253_/A1 _7277_/B _7253_/B _7952_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_171_383 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_171_372 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4465_ hold73/Z _4748_/I1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_117_28 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_89_117 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xhold368 _7575_/Q hold368/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
Xhold346 _7579_/Q hold346/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
Xhold357 hold357/I _7624_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
XFILLER_131_247 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6204_ hold47/Z _6208_/A2 _6204_/B _7737_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
Xhold379 _7898_/Q hold379/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
X_4396_ _7447_/Q input81/Z _4396_/S _4396_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_7184_ _7184_/A1 _7210_/A2 _7184_/B1 _7184_/B2 _7433_/Q _7185_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi221_1
X_6135_ hold406/Z _6140_/A2 _6136_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_98_673 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_640 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_651 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_6066_ hold41/Z _6072_/A2 _6066_/B hold439/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_112_494 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_97_172 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_662 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_673 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_684 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_695 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_5017_ _5230_/A1 _5024_/A2 _5200_/B _5529_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_4
XFILLER_172_9 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_38_250 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_38_272 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1806 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_66_592 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1839 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1828 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1817 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_81_584 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_81_551 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_26_69 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6968_ _7758_/Q _7202_/C2 _7201_/A2 _7748_/Q _6971_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_53_286 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_166_100 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5919_ hold90/Z hold276/I _5919_/B hold235/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_6899_ _7930_/Q _7133_/S _6900_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_167_667 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_22_673 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_42_46 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_182_604 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_139_369 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_108_734 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_150_534 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_122_247 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_3_29 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_1_577 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_49_537 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_49_548 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_76_367 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_76_356 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_64_518 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_57_570 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_17_489 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_44_242 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_60_735 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_9_611 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_158_656 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_157_122 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_157_144 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_8_132 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_172_103 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_8_176 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_160_309 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_148_90 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_126_531 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_153_383 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_113_225 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4250_ _7620_/Q _5954_/A1 _4812_/A1 _7494_/Q _4253_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_141_567 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4181_ _7733_/Q _6192_/A1 _4878_/A1 _7532_/Q _4868_/A1 _7528_/Q _4183_/A2 VDD VSS
+ gf180mcu_fd_sc_mcu7t5v0__aoi222_1
XFILLER_83_805 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_55_507 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_7940_ _7940_/D _7961_/RN _7940_/CLK _7940_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
X_7871_ _7871_/D _7961_/RN _7871_/CLK _7871_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffsnq_1
X_6822_ _7722_/Q _6881_/A2 _6881_/B1 _7698_/Q _6824_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_90_392 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_35_286 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6753_ _6753_/A1 _6753_/A2 _6753_/A3 _6754_/B2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor3_1
X_3965_ _7649_/Q _6005_/A1 _4231_/B1 input68/Z _3994_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_149_634 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3896_ _3896_/A1 _3896_/A2 _3896_/A3 _3918_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand3_2
X_5704_ _5704_/A1 _5704_/A2 _5704_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__and2_1
X_6684_ _6684_/A1 _6684_/A2 _6684_/A3 _6686_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor3_1
X_5635_ _5692_/B _5218_/C _5708_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_1
Xhold110 _7545_/Q _3643_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
X_5566_ _5602_/A2 _4993_/B _5663_/A1 _5566_/B _5567_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai31_1
X_5497_ _5452_/C _5498_/A2 _5497_/A3 _5499_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor3_1
Xhold121 _7339_/Q hold121/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
Xhold143 _7338_/Q hold143/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
X_4517_ hold47/Z _4521_/A2 _4517_/B hold545/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_7305_ input75/Z _4334_/Z _7305_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__and2_1
X_7236_ _3658_/I _7236_/A2 _7237_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_172_692 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_4448_ hold15/Z _4449_/A2 _4448_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__and2_4
XFILLER_132_534 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
Xhold154 _3793_/Z hold154/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
Xhold165 hold165/I hold165/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
XFILLER_104_247 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xhold176 hold176/I _5994_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
Xhold198 hold198/I _7422_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
XFILLER_144_37 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_104_258 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xhold187 _7896_/Q hold187/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
XFILLER_113_792 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_100_420 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_58_301 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_4379_ _4379_/I _7412_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_7167_ _7509_/Q _7191_/A2 _7190_/B1 _7468_/Q _7190_/A2 _7401_/Q _7168_/A2 VDD VSS
+ gf180mcu_fd_sc_mcu7t5v0__aoi222_1
X_7098_ _7779_/Q _7200_/A2 _7200_/B1 _7867_/Q _7100_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_6118_ hold433/Z _6123_/A2 _6119_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_86_676 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_492 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_481 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_470 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_46_507 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6049_ hold41/Z _6055_/A2 _6049_/B hold493/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_37_46 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_37_57 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_39_570 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2326 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2315 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2304 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2348 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2359 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2337 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1614 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1603 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_14_404 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1658 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1647 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1636 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1625 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_41_212 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1669 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_757 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_167_420 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_139_144 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_10_654 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
Xclkbuf_leaf_82_csclk clkbuf_leaf_9_csclk/I _7398_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_182_434 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_182_412 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_167_486 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_155_637 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_10_676 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_182_445 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_154_136 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_108_531 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_6_647 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_170_629 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_135_372 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xclkbuf_leaf_97_csclk _7558_/CLK _7561_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_123_578 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_123_567 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_78_53 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
Xclkbuf_leaf_20_csclk _7825_/CLK _7849_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_65_805 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_49_334 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_92_602 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_77_687 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_18_732 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
Xclkbuf_leaf_35_csclk clkbuf_3_7__f_csclk/Z _7755_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_17_231 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_150_80 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_72_392 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_17_275 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_17_286 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_18_798 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_32_212 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_177_228 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3750_ _7411_/Q _3774_/A2 _3751_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_158_453 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_173_434 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3681_ _7849_/Q _3681_/ZN VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_118_339 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_9_485 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5420_ _5062_/Z _5176_/B _5421_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_9_496 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_161_629 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_154_670 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xoutput215 _4410_/Z mgmt_gpio_out[15] VDD VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
Xoutput226 _7999_/Z mgmt_gpio_out[25] VDD VSS gf180mcu_fd_sc_mcu7t5v0__buf_8
X_5351_ _5498_/A2 _5622_/A1 _5534_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_114_501 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
Xoutput204 _3707_/ZN mgmt_gpio_oeb[5] VDD VSS gf180mcu_fd_sc_mcu7t5v0__buf_8
XFILLER_57_2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
Xoutput237 _4396_/Z mgmt_gpio_out[35] VDD VSS gf180mcu_fd_sc_mcu7t5v0__buf_8
X_4302_ _4308_/S _4296_/Z _7342_/Q _4303_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_114_534 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_99_223 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_99_212 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5282_ _5282_/A1 _5282_/A2 _5282_/A3 _5298_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand3_1
Xoutput259 _7568_/Q pll90_sel[2] VDD VSS gf180mcu_fd_sc_mcu7t5v0__buf_8
Xoutput248 _4436_/Z pad_flash_clk_oe VDD VSS gf180mcu_fd_sc_mcu7t5v0__buf_8
X_7021_ _7824_/Q _7202_/A2 _7204_/B1 _7768_/Q _7025_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_99_267 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_4233_ _7375_/Q hold114/I _6209_/A1 _7740_/Q _4256_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_114_29 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4164_ _7400_/Q _4589_/A1 _4527_/A1 _7374_/Q _4167_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_4095_ _7888_/Q _6520_/A1 _6209_/A1 _7742_/Q _4106_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_82_101 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_68_676 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_83_668 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_7923_ _7923_/D _7961_/RN _7938_/CLK _7923_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_67_197 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_55_326 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_55_337 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_70_318 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_70_307 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_24_713 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_36_540 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_169_707 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7854_ _7854_/D _7901_/RN _7881_/CLK _7854_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffsnq_1
XFILLER_63_370 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_23_212 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_23_223 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_24_735 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_169_718 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_169_729 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_168_206 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6805_ _7738_/Q _6878_/A2 _6805_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__or2_1
X_7785_ _7785_/D _7901_/RN _7865_/CLK _7785_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_51_543 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4997_ _3722_/I _3723_/I _5006_/B _5006_/C _5663_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand4_4
X_6736_ _7825_/Q _6891_/A2 _6891_/B1 _7671_/Q _6891_/C1 _7777_/Q _6738_/A3 VDD VSS
+ gf180mcu_fd_sc_mcu7t5v0__aoi222_1
XFILLER_176_250 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3948_ _3948_/A1 _3948_/A2 _3948_/A3 _3948_/A4 _3954_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand4_2
X_3879_ hold630/I _3869_/I hold55/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__or2_4
XFILLER_137_637 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6667_ _7684_/Q _6884_/B1 _6892_/B1 _7724_/Q _6681_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_5618_ _5689_/A1 _5692_/B _5618_/A3 _5618_/B1 _5620_/B _5632_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai32_1
X_6598_ _7434_/Q _7912_/Q _7911_/Q _6609_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_136_169 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_5549_ _5765_/A2 _5803_/A4 _5549_/A3 _5765_/A3 _5557_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand4_1
XFILLER_117_361 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_151_139 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_2_105 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xclkbuf_3_0__f_wb_clk_i clkbuf_0_wb_clk_i/Z _7912_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_160_673 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_144_191 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_105_567 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_78_407 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_78_429 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7219_ _7219_/A1 _7228_/S _7219_/B _7942_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_100_261 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_100_250 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_86_473 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_74_602 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2101 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_104_51 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_73_134 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_73_123 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_62_808 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2134 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2112 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2123 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_64_33 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2167 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2156 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_161_2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2145 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1433 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1422 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1411 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1400 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2189 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2178 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1455 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1466 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1444 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_64_99 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_15_779 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_42_554 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_54_392 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_159_228 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_120_72 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_1499 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1488 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1477 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_30_738 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_167_283 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_13_70 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_1_160 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_2_672 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_96_259 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_77_462 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_65_657 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_37_337 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_80_605 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_4920_ _4917_/Z _4919_/Z _4920_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__and2_4
XFILLER_18_584 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_52_318 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4851_ hold602/Z _4852_/A2 _4852_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_3802_ _7341_/Q _4383_/A1 _4306_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_21_716 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4782_ hold596/Z _4783_/A2 hold597/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_7570_ _7570_/D _7961_/RN _7570_/CLK _7570_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffsnq_2
XFILLER_158_250 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_146_412 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3733_ _4424_/A1 _3731_/Z _3733_/B _7980_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_6521_ hold750/Z _6536_/A2 _6522_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_173_242 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6452_ _6452_/A1 _7285_/A2 _6468_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_4
X_3664_ _3664_/I _4425_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__inv_1
X_5403_ _5579_/B _5591_/A2 _5559_/A1 _5577_/C _5407_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor4_1
XFILLER_134_629 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_173_286 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6383_ hold90/Z _6383_/A2 _6383_/B _7821_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_5334_ _5404_/A1 _5424_/A1 _5292_/B _5087_/B _5334_/C _5335_/A4 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi221_1
XFILLER_141_172 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_141_161 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_125_39 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_125_17 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5265_ _5624_/A1 _5759_/A1 _5724_/B _5561_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_87_215 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5196_ _5011_/B _3723_/I _5211_/A3 _4920_/Z _5209_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand4_2
X_7004_ _7702_/Q _7190_/C1 _7008_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_4216_ _3817_/I _4075_/B _4238_/B1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_96_771 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4147_ _4153_/A1 _4151_/A2 _4779_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_2
XFILLER_56_613 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_95_281 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_83_443 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_68_484 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_18_37 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4078_ _7670_/Q _6056_/A1 _5920_/A1 _7606_/Q _4219_/A2 input13/Z _4080_/A2 VDD VSS
+ gf180mcu_fd_sc_mcu7t5v0__aoi222_2
X_7906_ _7906_/D _7961_/RN _7940_/CLK _7906_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_2
X_7837_ _7837_/D _7901_/RN _7900_/CLK _7837_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_70_137 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_70_159 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_36_392 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_169_559 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_169_548 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_24_587 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7768_ _7768_/D _7901_/RN _7873_/CLK _7768_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffsnq_1
XFILLER_11_237 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_11_215 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_51_384 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_177_570 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_109_114 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7699_ _7699_/D _7961_/RN _7707_/CLK _7699_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
X_6719_ _7614_/Q _6647_/Z _6890_/A2 _7638_/Q _6720_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_7_219 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_149_283 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_137_445 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_20_782 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_137_489 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_3_425 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_3_469 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_133_684 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_132_172 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_182_78 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_120_345 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_59_440 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_120_389 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_115_61 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_87_760 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_101_570 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_46_112 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_47_624 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_62_605 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_46_156 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_47_668 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_34_318 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_34_329 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_131_93 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_91_20 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1241 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1230 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1274 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1263 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1252 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_70_671 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1296 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1285 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_7_775 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xhold709 _7373_/Q hold709/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
XFILLER_171_735 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_170_201 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_155_286 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_124_673 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_69_215 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5050_ _5006_/C _5448_/A1 _5179_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__and2_4
XFILLER_78_782 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_38_602 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4001_ _7552_/Q _4284_/A1 _4427_/B _4002_/B2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_93_774 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_1_73 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_38_668 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5952_ hold351/Z _5953_/A2 _5953_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_37_189 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_53_638 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4903_ _3723_/I _4946_/A1 _5648_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_4
XFILLER_18_392 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_178_334 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5883_ _4448_/Z _5885_/A2 _5883_/B _7586_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_33_340 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7622_ _7622_/D _7961_/RN _7643_/CLK _7622_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffsnq_1
X_4834_ hold621/Z _4835_/A2 hold622/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_178_389 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_166_529 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_159_570 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4765_ hold670/Z _4768_/A2 _4766_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_7553_ _7553_/D _7312_/Z _7977_/CLK _7553_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffnrnq_1
X_6504_ hold734/Z _6519_/A2 _6505_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_3716_ _7467_/Q _7210_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_147_776 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4696_ _3819_/Z _4460_/Z _4697_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_7484_ _7484_/D _7944_/CLK _7484_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_3647_ _7511_/Q _7214_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_161_212 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6435_ _6435_/A1 hold32/Z _6451_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_4
XFILLER_20_49 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6366_ hold90/Z _6366_/A2 _6366_/B _7813_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_115_651 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5317_ _5768_/A2 _5237_/Z _5624_/B _5648_/B2 _5326_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_1
Xhold14 hold14/I hold14/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
X_6297_ hold410/Z _6298_/A2 _6298_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_88_557 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
Xhold47 hold47/I hold47/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
Xhold36 hold36/I hold36/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
XFILLER_152_37 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5248_ _5338_/A1 _5369_/B _5303_/A3 _5618_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand3_2
XFILLER_130_676 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
Xhold25 hold25/I hold25/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
XFILLER_29_69 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
Xhold69 hold69/I hold69/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
Xhold58 hold58/I hold58/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
X_5179_ _5608_/B _5752_/B1 _5793_/A2 _5179_/B _5188_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai31_1
XFILLER_102_389 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_68_270 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_28_112 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_28_101 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_29_679 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_44_605 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_16_318 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_16_329 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_43_148 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_324 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_313 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_302 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_357 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_346 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_335 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_24_384 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_138_754 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_124_2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_137_286 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_153_779 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_4_756 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_106_673 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_105_150 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_126_93 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_35_638 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_34_148 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_62_479 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_15_351 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1082 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1071 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1060 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_15_373 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_30_310 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_30_321 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1093 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_156_540 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4550_ hold660/Z _4553_/A2 _4551_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_4481_ hold68/Z _4740_/I1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_143_212 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xhold506 _7892_/Q hold506/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
Xhold517 _7648_/Q hold517/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
X_6220_ hold269/Z _6225_/A2 hold270/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_144_757 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
Xhold528 hold528/I _7623_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
Xhold539 _7360_/Q hold539/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
X_6151_ hold41/Z _6157_/A2 _6151_/B _7712_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
XTAP_800 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_5102_ _5669_/A1 _5648_/A2 _5102_/B1 _5777_/A2 _5105_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XTAP_811 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_822 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_833 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_844 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_112_676 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_97_354 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6082_ hold507/Z _6089_/A2 _6083_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_855 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_866 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_877 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_5033_ _5199_/B _5201_/B _5369_/B _4944_/Z _5035_/A4 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor4_4
XFILLER_111_186 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_888 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_899 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_122_29 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_26_605 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_53_424 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6984_ _7847_/Q _7193_/A2 _7193_/B1 _7629_/Q _7193_/C1 _7725_/Q _6986_/A1 VDD VSS
+ gf180mcu_fd_sc_mcu7t5v0__aoi222_1
X_5935_ hold342/Z _5936_/A2 _5936_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_80_276 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_34_660 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_61_490 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5866_ hold68/Z _5868_/A2 _5866_/B _7579_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_34_682 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4817_ _7514_/Q _7959_/RN _4828_/S VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_4
XFILLER_21_354 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7605_ _7605_/D _7961_/RN _7648_/CLK _7605_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_166_337 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5797_ _5797_/A1 _5797_/A2 _5797_/B _5797_/C _5798_/A4 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XFILLER_181_318 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4748_ hold634/Z _4748_/I1 _4753_/S _7461_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_147_540 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_5_509 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_7536_ _7536_/D _7901_/RN _7895_/CLK _7536_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_174_392 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4679_ hold55/Z hold68/Z _4680_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_134_223 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_134_201 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_119_286 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7467_ _7467_/D _7961_/RN _7573_/CLK _7467_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
X_6418_ _6418_/A1 _7285_/A2 _6434_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_4
XFILLER_150_738 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_134_278 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_7398_ _7398_/D _7961_/RN _7398_/CLK _7398_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
X_6349_ hold90/Z _6349_/A2 _6349_/B _7805_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_115_481 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_88_321 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xinput115 wb_adr_i[28] _4368_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
Xinput104 wb_adr_i[18] _4924_/A4 VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
Xinput126 wb_adr_i[9] _4925_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_247 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xinput148 wb_dat_i[28] _7260_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
Xinput137 wb_dat_i[18] _7250_/B1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
Xinput159 wb_dat_i[9] _7245_/B1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_29_454 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_72_744 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_72_33 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_13_811 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_44_479 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_143 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_132 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_121 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_12_321 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_25_682 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_110 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_176 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_165 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_154 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_198 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_187 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_172_318 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_165_370 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_4_531 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_106_492 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_4_597 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_79_354 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_39_207 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_153_80 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_48_763 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_35_413 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_90_530 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3981_ _3981_/A1 _3981_/A2 _3981_/A3 _3990_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_90_552 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
X_5720_ hold23/I _5520_/C _5738_/C VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_16_671 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_31_641 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5651_ _5651_/A1 _5503_/C _5651_/A3 _5651_/A4 _5651_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__and4_1
XFILLER_87_2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_30_140 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5582_ _5578_/Z _5710_/A1 _5582_/A3 _5582_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__and3_1
XFILLER_129_551 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_117_702 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_30_195 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4602_ hold569/Z _4603_/A2 _4603_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_7321_ _7901_/RN _4334_/Z _7321_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_163_318 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_156_370 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4533_ hold676/Z _4548_/A2 _4534_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_7252_ _7252_/A1 _7280_/A2 _7277_/B _7252_/C _7253_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi211_1
Xhold303 _7751_/Q hold303/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
XFILLER_171_340 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_156_392 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
Xhold314 _3810_/S _3801_/S VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
Xhold325 _7768_/Q hold325/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
X_4464_ _7968_/Q _7506_/Q hold72/Z hold73/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_4
XFILLER_131_215 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_6203_ hold414/Z _6208_/A2 _6204_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
Xhold336 _7651_/Q hold336/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
Xhold369 _7786_/Q hold369/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
Xhold347 _7626_/Q hold347/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
Xhold358 _7874_/Q hold358/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
XFILLER_89_129 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_4395_ _7445_/Q input78/Z _4396_/S _4395_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_7183_ _7210_/A2 _7183_/A2 _7183_/A3 _7184_/B2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor3_1
XFILLER_140_760 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_100_602 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_98_685 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_6134_ hold41/Z _6140_/A2 _6134_/B _7704_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
XTAP_630 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_641 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_652 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_6065_ hold438/Z _6072_/A2 _6066_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_663 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_674 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_685 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_5016_ _5016_/A1 _5016_/A2 _5016_/B _5452_/C VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_4
XFILLER_85_357 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_696 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_26_413 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1807 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_26_37 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_54_744 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1829 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1818 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_81_563 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6967_ _6967_/A1 _6967_/A2 _6967_/A3 _6977_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_54_788 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5918_ hold234/Z hold276/I _5919_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_179_473 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_167_613 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6898_ _7433_/Q _7929_/Q _6898_/B1 _6898_/B2 _6900_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_167_657 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_167_635 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_22_663 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5849_ _7961_/RN _5849_/A2 _7285_/A2 _5851_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand3_1
X_7519_ _7519_/D _7959_/RN _7958_/CLK _7519_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_4
XFILLER_154_318 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_108_724 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_181_159 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_174_46 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_89_641 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_107_73 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_103_440 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_1_567 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_107_95 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_91_327 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_72_574 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_17_479 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_44_254 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_44_265 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_60_747 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_16_70 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_158_602 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_13_641 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_158_646 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_157_101 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_80_9 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_13_696 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_40_460 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_173_627 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_138_392 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_113_215 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_95_600 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4180_ _7685_/Q _6090_/A1 _4883_/A1 _7534_/Q _4893_/A1 _7538_/Q _4183_/A1 VDD VSS
+ gf180mcu_fd_sc_mcu7t5v0__aoi222_1
XFILLER_94_110 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_67_357 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_67_346 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_94_176 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_82_316 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7870_ _7870_/D _7961_/RN _7871_/CLK _7870_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffsnq_1
XFILLER_35_221 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6821_ _7658_/Q _6882_/B1 _6647_/Z _7618_/Q _6824_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_90_382 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_51_736 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6752_ _6752_/A1 _6752_/A2 _6752_/A3 _6752_/A4 _6753_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand4_1
X_3964_ hold25/Z hold156/Z _5828_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_4
X_5703_ _5104_/B _5658_/B _5685_/B _5247_/B _5703_/C _5704_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi221_1
X_6683_ _6683_/A1 _6683_/A2 _6683_/A3 _6683_/A4 _6684_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand4_1
X_3895_ input33/Z _4249_/A2 _4219_/A2 input19/Z _3896_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_2
XFILLER_176_443 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_164_605 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_5634_ _5790_/A1 _5726_/A1 _5634_/A3 _5634_/A4 _5637_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor4_1
XFILLER_136_329 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_136_318 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_128_17 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xhold100 _7450_/Q hold100/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
X_5565_ _5565_/A1 _5565_/A2 _5565_/A3 _5565_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__or3_1
XFILLER_163_137 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_129_381 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7304_ input75/Z _4334_/Z _7304_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__and2_1
Xhold144 _3785_/Z hold144/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
Xhold122 _3781_/Z hold122/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
XFILLER_132_513 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
Xhold111 hold111/I _3800_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
X_5496_ _5496_/A1 _4993_/B _5647_/A2 _5496_/B _5506_/C VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai31_1
Xhold133 hold133/I hold133/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
X_4516_ hold543/Z _4521_/A2 hold544/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_7235_ _7519_/Q _7235_/A2 _7238_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_4447_ input58/Z _3801_/S _4449_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
Xhold166 hold166/I _7436_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
XFILLER_104_237 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
Xhold177 hold177/I _7638_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
XFILLER_144_16 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
Xhold199 _7686_/Q hold199/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
Xhold188 hold188/I _7896_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
X_7166_ _7166_/A1 _7166_/A2 _7166_/A3 _7183_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_98_460 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6117_ hold41/Z _6123_/A2 _6117_/B _7696_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
Xclkbuf_leaf_1_csclk clkbuf_leaf_9_csclk/I _7589_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XTAP_460 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_4378_ _7964_/Q _4378_/A2 _7412_/Q _4379_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_7097_ _7097_/A1 _7097_/A2 _7097_/A3 _7097_/A4 _7106_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand4_1
XTAP_493 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_482 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_471 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_6048_ hold492/Z _6055_/A2 _6049_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_85_165 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_58_368 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_37_36 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2316 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2305 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_160_37 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_26_210 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_37_69 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_54_530 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2349 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2338 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2327 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1615 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1604 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1648 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1637 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1626 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_7999_ _7999_/I _7999_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_81_382 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_42_747 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1659 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_169_79 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_10_600 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_182_468 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_182_457 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_5_158 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_150_321 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_104_760 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_110_218 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_49_357 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_94_53 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_76_176 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_17_210 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_18_744 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_150_70 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_60_544 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_146_605 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_13_493 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_41_780 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_173_424 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_118_318 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3680_ _7857_/Q _3680_/ZN VDD VSS gf180mcu_fd_sc_mcu7t5v0__inv_1
XFILLER_9_475 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_145_148 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
Xoutput216 _7990_/Z mgmt_gpio_out[16] VDD VSS gf180mcu_fd_sc_mcu7t5v0__buf_8
X_5350_ _5689_/A2 _5687_/B _5350_/A3 _5788_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor3_1
Xoutput205 _3706_/ZN mgmt_gpio_oeb[6] VDD VSS gf180mcu_fd_sc_mcu7t5v0__buf_8
Xoutput238 _4387_/Z mgmt_gpio_out[36] VDD VSS gf180mcu_fd_sc_mcu7t5v0__buf_8
X_4301_ _4301_/A1 _4301_/A2 _7343_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
Xoutput227 _8000_/Z mgmt_gpio_out[26] VDD VSS gf180mcu_fd_sc_mcu7t5v0__buf_8
XFILLER_126_384 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_114_546 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5281_ _5685_/B _5292_/B _5585_/C _5282_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi21_1
Xoutput249 _4417_/Z pad_flash_csb VDD VSS gf180mcu_fd_sc_mcu7t5v0__buf_8
X_7020_ _7760_/Q _7202_/C2 _7202_/B1 _7784_/Q _7025_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_102_708 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4232_ input34/Z _4232_/A2 _4848_/A1 _7509_/Q _4260_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_4_62 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_110_741 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4163_ _7376_/Q hold114/I _6452_/A1 _7855_/Q _7584_/Q _5874_/A1 _4167_/A1 VDD VSS
+ gf180mcu_fd_sc_mcu7t5v0__aoi222_1
XFILLER_67_132 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4094_ _7760_/Q _6248_/A1 _5817_/A1 _7560_/Q _6333_/A1 _7800_/Q _4106_/A2 VDD VSS
+ gf180mcu_fd_sc_mcu7t5v0__aoi222_2
XFILLER_95_496 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_82_135 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_82_124 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7922_ _7922_/D _7961_/RN _7938_/CLK _7922_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
X_7853_ _7853_/D _7901_/RN _7853_/CLK _7853_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_82_179 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_4996_ _3722_/I _3723_/I _5006_/B _5006_/C _4996_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__and4_4
X_7784_ _7784_/D _7901_/RN _7899_/CLK _7784_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffsnq_1
X_6804_ _7133_/S _6804_/A2 _6804_/B _7926_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_24_747 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_51_555 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_149_421 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6735_ _7761_/Q _6892_/A2 _6893_/C1 _7631_/Q _6738_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_3947_ _7788_/Q _6299_/A1 _5988_/A1 _7642_/Q _3948_/A4 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_51_566 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_139_16 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_176_273 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3878_ hold630/I _3869_/I _4231_/B1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_4
X_6666_ _7668_/Q _6891_/B1 _6880_/B1 _7806_/Q _6677_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_136_126 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5617_ _5618_/B1 _5620_/B _5617_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__or2_1
X_6597_ _7912_/Q _7911_/Q _6953_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_4
X_5548_ _5548_/A1 _5548_/A2 _5548_/A3 _5765_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_132_321 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_105_524 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_160_663 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5479_ _5779_/A1 _5479_/A2 _5503_/C VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_7218_ _7942_/Q _7228_/S _7219_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_99_780 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7149_ _7699_/Q _7194_/A2 _7190_/B1 _7619_/Q _7153_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_171_69 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_101_774 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_86_463 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_58_165 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_58_198 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2135 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2113 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2124 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2102 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_73_157 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_64_45 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_27_552 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2168 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2157 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2146 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1423 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1412 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1401 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_511 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_54_371 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2179 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_154_2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1445 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1456 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1434 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_544 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_120_84 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1489 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1478 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1467 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_128_605 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_168_796 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_127_115 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_167_295 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_155_446 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_10_463 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_143_619 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_129_82 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_6_456 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_163_490 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_151_630 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_151_641 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_123_354 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_69_419 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_49_132 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_77_496 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_65_636 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_64_124 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_161_91 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_18_530 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_64_179 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_60_330 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4850_ _4448_/Z _4852_/A2 _4850_/B _7509_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_3801_ _3801_/I0 hold131/Z _3801_/S _3801_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_4
XTAP_1990 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_60_396 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4781_ _4448_/Z _4783_/A2 _4781_/B _7476_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_6520_ _6520_/A1 _7285_/A2 _6536_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_4
XFILLER_174_700 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_158_273 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_146_402 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_119_638 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3732_ _7965_/Q _3731_/Z _3733_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_174_744 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6451_ hold90/Z _6451_/A2 _6451_/B _7853_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_9_294 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_9_283 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3663_ _3663_/I _4392_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_5402_ _5689_/A1 _5405_/B _5504_/A3 _5372_/Z _5576_/B2 _5577_/C VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai32_1
XFILLER_146_479 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6382_ hold236/Z _6383_/A2 _6383_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_5333_ _5689_/A2 _5687_/B _5333_/A3 _5495_/B2 _5258_/B _5334_/C VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai32_1
XFILLER_114_321 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5264_ _5714_/B1 _5687_/B _5504_/A3 _5701_/C _5287_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai31_1
XFILLER_125_29 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_88_728 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5195_ _5087_/C _4914_/Z _5210_/A3 _5195_/B _5209_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai31_1
XFILLER_102_549 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4215_ _7980_/Q _7965_/Q _7573_/Q _4215_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__or3_1
X_7003_ _7003_/A1 _7133_/S _7003_/B1 _7003_/B2 _7932_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_110_560 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_68_463 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
Xclkbuf_leaf_81_csclk clkbuf_leaf_9_csclk/I _7802_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
X_4146_ _4153_/A1 _4155_/A2 _4769_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_2
XFILLER_95_293 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_28_316 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4077_ input45/Z _4275_/A2 _5937_/A1 _7614_/Q _7646_/Q _6005_/A1 _4080_/A1 VDD VSS
+ gf180mcu_fd_sc_mcu7t5v0__aoi222_2
XFILLER_83_488 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_83_499 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_70_105 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7905_ _7905_/D _7961_/RN _7940_/CLK _7905_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
X_7836_ _7836_/D _7901_/RN _7883_/CLK _7836_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
Xclkbuf_leaf_96_csclk _7558_/CLK _7565_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_34_37 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4979_ _5069_/A2 _4930_/Z _4979_/A3 _4953_/Z _5366_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand4_4
XFILLER_140_8 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7767_ _7767_/D _7901_/RN _7895_/CLK _7767_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffsnq_1
XFILLER_51_396 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7698_ _7698_/D _7961_/RN _7698_/CLK _7698_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
X_6718_ _7718_/Q _6881_/A2 _6885_/B1 _7710_/Q _6720_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_6649_ _7910_/Q _6658_/A2 _6658_/A3 _6890_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor3_4
XFILLER_180_747 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
Xclkbuf_leaf_34_csclk clkbuf_3_7__f_csclk/Z _7810_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_118_682 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_118_671 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_180_769 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_133_641 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_105_354 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_182_68 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
Xclkbuf_leaf_49_csclk clkbuf_3_6__f_csclk/Z _7691_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_115_73 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_115_51 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_87_772 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_87_783 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_74_400 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_59_496 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_19_327 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_46_102 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_75_66 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_75_77 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_131_50 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_61_116 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_46_179 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_1231 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1220 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_330 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_54_190 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_55_691 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1275 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1264 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1253 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1242 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_15_566 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1297 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1286 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_175_519 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
Xclkbuf_3_4__f_csclk clkbuf_0_csclk/Z _7592_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_30_569 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_156_744 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_156_733 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_11_783 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_10_260 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_6_264 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_170_257 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_41_6 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_124_685 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_85_709 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_111_357 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4000_ _4206_/A1 _7227_/I0 _4002_/B1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_1_30 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_65_455 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_37_157 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_5951_ hold68/Z _5953_/A2 _5951_/B hold403/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_65_499 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_52_105 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_52_116 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4902_ _5309_/A1 _3723_/I _5666_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_61_661 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_61_650 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5882_ hold712/Z _5885_/A2 _5883_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_7621_ _7621_/D _7961_/RN _7627_/CLK _7621_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffsnq_1
X_4833_ _4448_/Z _4835_/A2 _4833_/B _7504_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_178_379 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_147_722 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_147_700 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4764_ _4764_/A1 _7285_/A2 _4768_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_7552_ _7552_/D _7311_/Z _7977_/CLK _7552_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffnrnq_1
XFILLER_174_530 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_146_210 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6503_ _6503_/A1 _7285_/A2 _6519_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_4
X_7483_ _7483_/D _7944_/CLK _7483_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_3715_ _7466_/Q _7184_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_146_265 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_146_254 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4695_ hold170/Z _4718_/A1 _4698_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_6434_ hold90/Z _6434_/A2 _6434_/B _7845_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_3646_ _7516_/Q _5678_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__inv_1
XFILLER_162_747 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_161_202 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_147_799 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6365_ hold230/Z _6366_/A2 _6366_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_115_641 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6296_ hold68/Z _6298_/A2 _6296_/B _7780_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_130_600 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5316_ _5685_/B _5648_/B2 _5316_/B _5316_/C _5356_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XFILLER_114_162 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_130_655 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_102_346 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5247_ _5685_/B _5724_/B _5247_/B _5288_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_88_547 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xhold37 hold37/I hold37/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
Xhold15 hold15/I hold15/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
XFILLER_69_761 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xhold26 hold26/I hold26/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
Xhold48 hold48/I hold48/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
X_5178_ _5178_/A1 _5178_/A2 _5178_/A3 _5188_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor3_1
Xhold59 hold59/I hold59/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
XFILLER_69_783 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_56_411 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_4129_ _4217_/A2 hold25/Z _4759_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_28_179 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_83_296 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_24_330 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_325 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_314 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_303 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_40_812 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_358 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_347 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_169_357 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_336 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
X_7819_ _7819_/D _7901_/RN _7819_/CLK _7819_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_101_53 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_138_700 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_101_97 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_61_46 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_138_744 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_137_210 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_137_232 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_152_202 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_117_2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_180_555 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_180_544 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_4_768 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_3_212 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_180_599 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_161_780 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_121_633 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_79_547 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_121_655 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_86_32 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_67_709 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_121_699 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_120_198 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_120_176 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_87_580 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_47_411 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_19_70 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_47_444 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_90_723 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_34_105 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_47_499 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_34_116 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_31_812 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_43_672 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1083 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1072 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1061 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1050 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_89_6 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1094 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_128_254 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4480_ _7971_/Q _7506_/Q hold67/Z hold68/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_4
XFILLER_171_511 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_156_596 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_144_747 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_116_438 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
Xhold507 _7680_/Q hold507/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
Xhold518 hold518/I _7648_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
XFILLER_171_566 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_171_555 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_144_769 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_143_224 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_116_449 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
Xhold529 _7873_/Q hold529/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
X_6150_ hold291/Z _6157_/A2 _6151_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_124_460 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_98_812 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_801 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_151_290 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5101_ _5602_/A1 _5647_/A2 _5777_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_2
XFILLER_32_2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_812 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_823 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_834 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_6081_ hold73/Z _6089_/A2 _6081_/B _7679_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
XTAP_845 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_856 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_867 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_57_208 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5032_ _4965_/B _5366_/A2 _5608_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_4
XFILLER_111_176 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_78_580 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_878 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_889 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_38_433 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_81_712 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_38_488 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6983_ _7677_/Q _7191_/A2 _7191_/B1 _7799_/Q _6992_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_53_436 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5934_ hold68/Z _5936_/A2 _5934_/B _7610_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_81_789 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_80_266 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_40_108 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_53_469 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_5865_ hold346/Z _5868_/A2 _5866_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_22_812 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_33_171 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_34_672 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_178_176 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_166_316 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4816_ _4454_/Z _4816_/A2 _4816_/B hold588/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_7604_ _7604_/D _7961_/RN _7645_/CLK _7604_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffsnq_1
XFILLER_21_344 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5796_ _5785_/B _5795_/Z _5806_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_4747_ hold9/Z hold7/Z _4753_/S hold10/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_7535_ _7535_/D _7901_/RN _7895_/CLK _7535_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_174_382 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_162_500 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_4678_ _7430_/Q _4685_/A1 _4681_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_107_438 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_7466_ _7466_/D _7961_/RN _7573_/CLK _7466_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
X_6417_ hold90/Z _6417_/A2 _6417_/B _7837_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_7397_ _7397_/D _7961_/RN _7874_/CLK _7397_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_150_717 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_134_268 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6348_ hold376/Z _6349_/A2 _6349_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_89_812 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_143_780 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_115_493 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_1_749 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
Xinput127 wb_cyc_i _4366_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
Xinput116 wb_adr_i[29] _4372_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
Xinput105 wb_adr_i[19] _4924_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_130_463 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_6279_ hold68/Z _6281_/A2 _6279_/B _7772_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_102_132 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xinput149 wb_dat_i[29] _7264_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
Xinput138 wb_dat_i[19] _7254_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_130_485 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_102_176 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_16_105 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_57_775 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_112_52 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_29_499 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_112_85 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_112_74 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_32_609 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_44_458 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_100 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_169_110 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_133 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_122 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_111 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_166 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_155 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_144 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_199 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_188 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_177 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_173_809 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_126_747 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_4_521 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_180_352 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_153_566 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_106_460 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_98_108 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_133_290 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_79_344 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_153_70 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_121_496 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_67_517 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_760 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_39_219 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_94_358 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_48_731 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_48_753 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_75_550 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_75_561 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_63_712 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_35_425 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3980_ _7681_/Q _6073_/A1 hold119/I _7729_/Q _3981_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_63_778 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_62_266 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_35_469 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_15_160 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_22_108 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_50_439 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_5650_ _3728_/I _5122_/Z _5650_/A3 _5651_/A4 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_176_647 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_4601_ _4448_/Z _4603_/A2 _4601_/B _7403_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_164_809 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5581_ _5212_/Z _5702_/A2 _5581_/B _5581_/C _5582_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XFILLER_129_541 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7320_ _7901_/RN _4334_/Z _7320_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__and2_1
X_4532_ hold114/Z hold32/Z _4548_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_4
XFILLER_116_213 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_116_202 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_7_73 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_7251_ _7251_/A1 _7251_/A2 _7252_/C VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_4463_ _7506_/Q _7258_/A1 hold72/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
Xhold315 _7794_/Q hold315/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
Xhold304 _7795_/Q hold304/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
Xhold326 _7880_/Q hold326/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
XFILLER_171_352 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6202_ hold41/Z _6208_/A2 _6202_/B _7736_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
Xhold337 hold337/I _7651_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
Xhold348 hold348/I _7626_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
Xhold359 _7625_/Q hold359/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
XFILLER_125_780 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4394_ _7444_/Q input80/Z _4396_/S _4394_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_7182_ _7182_/A1 _7182_/A2 _7182_/A3 _7183_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_86_804 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6133_ hold451/Z _6140_/A2 _6134_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_620 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_631 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_642 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_133_29 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_112_496 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_112_463 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_6064_ hold73/Z _6072_/A2 _6064_/B hold425/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
XTAP_653 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_664 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_675 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_686 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_5015_ _5139_/A1 _5014_/Z _5015_/B _5538_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi21_4
XTAP_697 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1819 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1808 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_81_553 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6966_ _7790_/Q _7190_/A2 _7194_/C1 _7806_/Q _6966_/C _6967_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi221_1
XFILLER_26_458 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5917_ hold68/Z hold276/Z _5917_/B _7602_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_81_586 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_41_428 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6897_ _7210_/A1 _6767_/C _7433_/Q _6898_/B2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_179_496 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5848_ _4448_/Z _5848_/A2 _5848_/B hold755/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_21_141 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_42_37 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_158_37 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5779_ _5779_/A1 _5779_/A2 _5779_/B1 _5292_/B _5780_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_182_639 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_182_628 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_166_179 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_7518_ _7518_/D _7959_/RN _7958_/CLK _7518_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_4
XFILLER_108_747 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_162_352 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_150_514 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_7449_ _7449_/D input75/Z _7865_/CLK _7449_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_103_430 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_1_557 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_131_783 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_1_579 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_130_282 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_103_496 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_88_196 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_67_67 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_76_369 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_45_712 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_123_73 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_83_33 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_72_531 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_17_425 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_29_296 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_17_469 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_25_491 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_172_105 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_32_92 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_32_81 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_172_138 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_148_92 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_107_791 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_99_428 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_79_141 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_94_133 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_94_144 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_94_122 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_94_155 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_63_531 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_6820_ _7650_/Q _6880_/C2 _6892_/A2 _7764_/Q _6824_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_23_428 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_35_288 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6751_ _7663_/Q _6885_/A2 _6885_/B1 _7711_/Q _6752_/A4 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_3963_ hold19/Z _3787_/Z hold127/Z _3963_/A4 _3963_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__or4_4
XFILLER_50_247 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_176_433 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5702_ _5212_/Z _5702_/A2 _5702_/B _5702_/C _5782_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi211_2
X_3894_ _7805_/Q _6333_/A1 _5988_/A1 _7643_/Q _3896_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_6682_ _7798_/Q _6883_/A2 _6890_/B1 _7846_/Q _6683_/A4 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_5633_ _5614_/Z _5622_/Z _5684_/A2 _5633_/A4 _5634_/A4 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand4_1
X_5564_ _5565_/A1 _5565_/A2 _5565_/A3 _5578_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor3_1
XFILLER_148_179 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_129_371 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_12_29 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xhold101 hold101/I hold101/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
XFILLER_157_691 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_4515_ hold41/Z _4521_/A2 _4515_/B hold553/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_7303_ input75/Z _4334_/Z _7303_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_160_812 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5495_ _4993_/B _5647_/A2 _5797_/A2 _5687_/C _5495_/B2 _5742_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai32_1
Xhold123 hold123/I hold123/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
XFILLER_105_706 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xhold134 hold134/I hold134/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
X_7234_ _3658_/I _7281_/C2 _7235_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_4446_ _7506_/Q hold14/Z hold15/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
Xhold167 _7599_/Q hold167/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
XFILLER_104_227 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_104_205 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xhold156 _3963_/Z hold156/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
Xhold189 _7888_/Q hold189/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
Xhold178 _7856_/Q hold178/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
X_4377_ _7965_/Q _4327_/S _4378_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_7165_ _7373_/Q _7203_/B1 _7204_/A2 _7399_/Q _7166_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_113_783 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6116_ hold452/Z _6123_/A2 _6117_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_450 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_7096_ _7380_/Q _7188_/A2 _7096_/B _7097_/A4 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_58_336 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_58_325 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_494 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_483 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_461 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_472 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_6047_ hold73/Z _6055_/A2 _6047_/B hold294/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_100_455 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_85_144 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_27_701 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_27_712 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_37_48 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2317 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2306 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_37_59 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2339 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2328 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1605 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_27_767 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1649 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1638 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1627 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1616 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_7998_ _7998_/I _7998_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_14_406 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_26_266 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_27_789 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_42_726 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6949_ _6949_/I _7210_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_3
XFILLER_169_58 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_22_472 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_167_499 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_154_105 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_139_168 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_6_605 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_123_503 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_78_33 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_2_811 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
Xhold690 _7376_/Q hold690/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
XFILLER_89_461 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_1_354 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_77_645 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_77_689 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_92_637 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_27_70 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_33_704 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_150_60 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_72_372 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_60_501 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_45_597 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_60_534 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_32_247 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_41_792 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_145_116 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_71_6 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_145_127 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
Xoutput217 _7991_/Z mgmt_gpio_out[17] VDD VSS gf180mcu_fd_sc_mcu7t5v0__buf_8
XFILLER_160_108 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_142_812 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_126_330 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xoutput206 _3705_/ZN mgmt_gpio_oeb[7] VDD VSS gf180mcu_fd_sc_mcu7t5v0__buf_8
Xoutput239 _4386_/Z mgmt_gpio_out[37] VDD VSS gf180mcu_fd_sc_mcu7t5v0__buf_8
X_4300_ _3812_/Z _4297_/Z _4300_/B _4300_/C _4301_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai211_1
Xoutput228 _8001_/Z mgmt_gpio_out[27] VDD VSS gf180mcu_fd_sc_mcu7t5v0__buf_8
X_5280_ _5482_/B2 _5292_/B _5690_/A1 _5575_/A2 _5412_/B _5282_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi221_1
X_4231_ input71/Z _5903_/A1 _4231_/B1 input36/Z _4280_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_141_366 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_4162_ _4162_/A1 _4162_/A2 _4162_/A3 _4204_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand3_2
XFILLER_110_764 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_4093_ _7816_/Q hold134/I _6316_/A1 _7792_/Q hold26/I _7577_/Q _4106_/A1 VDD VSS
+ gf180mcu_fd_sc_mcu7t5v0__aoi222_2
XFILLER_83_604 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_67_144 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_83_637 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_67_199 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7921_ _7921_/D _7961_/RN _7938_/CLK _7921_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_55_339 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_70_309 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_36_531 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7852_ _7852_/D _7901_/RN _7852_/CLK _7852_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_63_361 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_63_372 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_51_523 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_169_709 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4995_ _5602_/A2 _4993_/B _4993_/C _4998_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor3_1
X_6803_ _7926_/Q _7133_/S _6804_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_7783_ _7783_/D _7901_/RN _7887_/CLK _7783_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffsnq_1
XFILLER_51_545 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6734_ _7727_/Q _6892_/B1 _6738_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_3946_ _7618_/Q _5937_/A1 _6226_/A1 _7754_/Q _7804_/Q _6333_/A1 _3948_/A3 VDD VSS
+ gf180mcu_fd_sc_mcu7t5v0__aoi222_2
XFILLER_23_28 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_136_105 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3877_ _4153_/A1 hold128/Z _6005_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_4
X_6665_ _7910_/Q _6665_/A2 _6665_/A3 _6665_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__and3_2
XFILLER_149_499 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5616_ _5616_/A1 _5643_/B1 _5176_/B _5620_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor3_4
X_6596_ _7434_/Q _6599_/A2 _6596_/B _7911_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_5547_ _5547_/A1 _5547_/A2 _5764_/A2 _5646_/A2 _5549_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor4_1
XFILLER_133_812 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5478_ _5797_/A1 _5543_/C _5543_/B _5545_/B _5662_/A1 _5505_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai32_1
X_7217_ _7517_/D _7959_/RN _7228_/S VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_4
X_4429_ _4400_/S input68/Z _4429_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_113_580 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_7148_ _7148_/A1 _7148_/A2 _7148_/A3 _7159_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_58_133 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_101_764 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_100_252 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7079_ _7079_/A1 _7210_/A2 _7433_/Q _7080_/B2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_74_615 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_47_807 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_100_263 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_74_637 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2114 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2125 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2103 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_27_542 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2158 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2147 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2136 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1424 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1413 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1402 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_54_361 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2169 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1446 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1457 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1435 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_14_247 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_42_534 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_147_2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_120_52 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1479 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1468 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_80_34 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_127_105 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_10_453 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_155_425 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_182_244 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_142_108 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_89_21 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_163_480 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_124_812 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_108_396 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_97_707 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_151_686 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_49_144 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_92_434 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_64_103 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_49_177 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_38_91 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_80_629 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_61_810 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_73_692 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_72_191 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3800_ _7506_/Q hold131/Z _3800_/B _3850_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_4
X_4780_ hold651/Z _4783_/A2 _4781_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_159_753 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_1991 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1980 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_60_375 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3731_ _3744_/A1 _7411_/Q _3730_/Z _3731_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__and3_1
Xclkbuf_leaf_0_csclk clkbuf_leaf_9_csclk/I _7886_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
X_6450_ hold409/Z _6451_/A2 _6451_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_3662_ _7415_/Q _4380_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_6381_ hold68/Z _6383_/A2 _6381_/B _7820_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_5401_ _5673_/A1 _5706_/A2 _5401_/A3 _5401_/A4 _5414_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand4_1
XFILLER_62_2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_161_428 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5332_ _5258_/B _5495_/B2 _5757_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_115_812 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_141_141 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5263_ _5433_/C _5768_/A3 _5681_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_88_718 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_87_217 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5194_ _5199_/B _3727_/I _4915_/Z _4996_/Z _5371_/C VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand4_4
XFILLER_87_239 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4214_ hold20/Z _4075_/B hold21/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_7002_ _7931_/Q _6556_/B _7002_/B _7003_/B2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_68_442 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4145_ _4153_/A1 _3869_/I _4843_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_95_283 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_83_423 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_83_412 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_141_29 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4076_ _7880_/Q _6503_/A1 _4104_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_83_467 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_70_117 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7904_ _7904_/D _7961_/RN _7940_/CLK _7904_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_52_810 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7835_ _7835_/D _7901_/RN _7883_/CLK _7835_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_64_692 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_24_534 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4978_ _5104_/B _5669_/B _4999_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_7766_ _7766_/D _7901_/RN _7881_/CLK _7766_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffsnq_1
XFILLER_165_712 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_137_414 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_7697_ _7697_/D _7961_/RN _7707_/CLK _7697_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
X_6717_ _7646_/Q _6880_/C2 _6882_/B1 _7654_/Q _6720_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_3929_ hold124/I _4075_/B _4176_/C VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_2
XFILLER_177_583 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_164_211 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_149_274 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_109_127 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6648_ _6878_/A2 _6663_/A4 _6664_/A2 _6880_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor3_4
XFILLER_50_37 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_166_37 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_124_108 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_117_171 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_117_160 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_106_812 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6579_ _7907_/Q _7906_/Q _6663_/A4 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_4
XFILLER_59_57 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_59_46 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_115_41 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_86_250 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_87_795 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_46_114 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_47_626 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_86_294 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_61_106 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_131_73 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_1232 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1221 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1210 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_27_394 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_131_95 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1265 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1254 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1243 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_70_673 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_30_504 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1298 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1287 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1276 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_30_515 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_168_550 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_10_250 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_128_458 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_143_428 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_7_799 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_170_247 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_123_130 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_2_460 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_93_721 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_77_283 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_65_423 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_65_412 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_92_242 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5950_ hold402/Z _5953_/A2 _5951_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_4901_ _3722_/I _5006_/B _5006_/C _4946_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand3_4
XFILLER_80_448 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_7620_ _7620_/D _7961_/RN _7627_/CLK _7620_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffsnq_1
X_5881_ _5881_/A1 _7285_/A2 _5885_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_60_183 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4832_ hold710/Z _4835_/A2 _4833_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_147_712 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_4763_ _4454_/Z _4763_/A2 _4763_/B _7469_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_7551_ _7551_/D _7310_/Z _4418_/I1 _7551_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffnrnq_1
XFILLER_119_425 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4694_ _4718_/A1 hold162/Z _4694_/B hold163/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_6502_ hold90/Z _6502_/A2 _6502_/B _7877_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_3714_ _7611_/Q _6849_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_7482_ _7482_/D _7949_/CLK _7482_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_147_767 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_119_469 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6433_ hold463/Z _6434_/A2 _6434_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_174_575 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_3645_ _7517_/Q _4376_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_106_108 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_20_29 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_161_247 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6364_ hold68/Z _6366_/A2 _6364_/B _7812_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_136_29 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5315_ _5545_/A2 _5687_/B _5648_/B2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_4
X_6295_ hold449/Z _6298_/A2 _6296_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_419 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5246_ _5199_/B _5201_/B _5421_/A1 _5333_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_114_174 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
Xhold38 hold38/I hold38/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
Xhold16 hold16/I hold16/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
Xhold27 hold27/I hold27/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
XFILLER_29_49 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
Xhold49 hold49/I hold49/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
X_5177_ _5651_/A1 _5769_/A1 _5177_/A3 _5178_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_68_250 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4128_ hold118/Z _4151_/A2 _4868_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_4059_ _7849_/Q _6435_/A1 _6265_/A1 _7769_/Q _4232_/A2 input6/Z _4063_/A1 VDD VSS
+ gf180mcu_fd_sc_mcu7t5v0__aoi222_1
XFILLER_16_309 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_83_286 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_315 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_304 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_359 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_348 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_169_347 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_337 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_326 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
X_7818_ _7818_/D _7901_/RN _7818_/CLK _7818_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_24_375 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_52_673 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7749_ _7749_/D _7901_/RN _7753_/CLK _7749_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffsnq_1
XFILLER_137_222 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_125_428 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_180_534 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_152_247 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_137_299 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_4_747 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_105_130 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_79_515 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_106_697 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_120_144 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_94_529 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_87_570 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_47_423 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_19_82 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_142_61 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_90_713 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_16_810 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_47_478 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_62_459 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1040 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1073 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1062 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1051 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_35_92 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_42_172 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_175_317 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_129_712 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_1095 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1084 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_156_531 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_30_389 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_11_570 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
Xhold508 _7836_/Q hold508/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
XFILLER_143_236 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
Xhold519 _7843_/Q hold519/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
XFILLER_98_802 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xclkbuf_leaf_95_csclk _7558_/CLK _7567_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
X_5100_ _5705_/A2 _5585_/A1 _5573_/C _5105_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_6080_ hold445/Z _6089_/A2 _6081_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_802 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_813 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_824 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_835 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_111_144 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_111_133 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_5031_ _5104_/B _5658_/B _5031_/B _5038_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_97_345 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_846 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_857 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_868 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_112_689 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_85_518 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_25_2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_879 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_66_743 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_66_798 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_25_106 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_38_478 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_65_286 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_6982_ _7791_/Q _7190_/A2 _7190_/B1 _7613_/Q _7190_/C1 _7701_/Q _6992_/A2 VDD VSS
+ gf180mcu_fd_sc_mcu7t5v0__aoi222_1
XFILLER_53_448 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
Xclkbuf_leaf_33_csclk clkbuf_3_7__f_csclk/Z _7852_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
X_5933_ hold378/Z _5936_/A2 _5934_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_80_245 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5864_ hold47/Z _5868_/A2 _5864_/B _7578_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_33_161 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7603_ _7603_/D _7901_/RN _7603_/CLK _7603_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
X_4815_ hold587/Z _4816_/A2 _4816_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_5795_ _5795_/A1 _5795_/A2 _5795_/A3 _5795_/A4 _5795_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__or4_1
X_7534_ _7534_/D _7961_/RN _7642_/CLK _7534_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
X_4746_ _4454_/Z _4753_/S _4746_/B _7459_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_147_542 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xclkbuf_leaf_48_csclk clkbuf_3_6__f_csclk/Z _7818_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
X_7465_ _7465_/D _7901_/RN _7583_/CLK _7465_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
X_4677_ _4685_/A1 hold49/Z _4677_/B hold50/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_147_39 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_107_428 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_162_534 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_135_759 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_134_247 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6416_ hold450/Z _6417_/A2 _6417_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_7396_ _7396_/D _7961_/RN _7396_/CLK _7396_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_134_258 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6347_ hold68/Z _6349_/A2 _6347_/B _7804_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_122_409 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_103_601 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_1_706 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_102_100 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_216 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
Xinput117 wb_adr_i[2] _5006_/C VDD VSS gf180mcu_fd_sc_mcu7t5v0__buf_12
Xinput106 wb_adr_i[1] _3722_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__buf_12
X_6278_ hold461/Z _6281_/A2 _6279_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_102_144 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
Xinput139 wb_dat_i[1] _7247_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
Xinput128 wb_dat_i[0] _7242_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_102_166 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_5229_ _5290_/B _5645_/A3 _5573_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_88_389 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_69_570 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_69_592 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_56_69 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_57_765 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_112_42 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_112_31 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_112_20 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_71_212 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_72_57 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_134 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_123 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_12_312 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_101 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_112 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_169_166 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_169_144 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_167 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_156 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_145 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_189 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_178 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_40_676 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_138_531 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_12_389 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_8_338 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_138_575 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_125_203 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_141_707 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_140_206 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_134_770 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_180_397 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_97_54 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_153_60 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_121_486 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_121_475 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_772 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_153_93 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_47_286 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_16_651 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_50_407 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_16_673 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4600_ hold714/Z _4603_/A2 _4601_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_5580_ _5580_/A1 _5636_/A1 _5380_/I _5581_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__or3_1
X_4531_ _4454_/Z _4531_/A2 _4531_/B _7374_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_7250_ _7520_/Q _7250_/A2 _7250_/B1 _7518_/Q _7251_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_144_534 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_144_523 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
Xhold305 hold305/I _6328_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
Xhold316 _7840_/Q hold316/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
X_4462_ _4487_/A1 _4460_/Z _4462_/B hold248/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
Xhold327 _7720_/Q hold327/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
X_6201_ hold446/Z _6208_/A2 _6202_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_116_247 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xhold349 _7739_/Q hold349/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
Xhold338 _7659_/Q hold338/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
XFILLER_125_792 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4393_ _7881_/Q _4396_/S _4393_/B _4393_/ZN VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_2
X_7181_ _7371_/Q _7201_/A2 _7205_/B1 _7537_/Q _7182_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_140_751 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_112_431 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6132_ hold73/Z _6140_/A2 _6132_/B _7703_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_98_676 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_610 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_621 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_632 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_643 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_112_486 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_6063_ hold424/Z _6072_/A2 _6064_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_100_615 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_100_626 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_58_529 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_654 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_665 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_676 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_5014_ _5195_/B _4926_/Z _5010_/Z _5014_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__or3_2
XFILLER_100_637 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_85_337 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_687 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_698 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_26_404 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_39_765 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_39_776 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_93_392 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_81_510 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_66_584 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_53_201 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_1809 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_6965_ _6965_/A1 _6965_/A2 _6965_/A3 _6966_/C VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand3_1
X_5916_ hold85/Z hold276/I _5917_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_81_598 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_22_621 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6896_ _6888_/Z _6896_/A2 _6896_/A3 _6895_/Z _6898_/B1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand4_1
XFILLER_166_125 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5847_ _7571_/Q _5848_/A2 _5848_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_22_676 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5778_ _5778_/A1 _5737_/B _5710_/Z _5733_/Z _5785_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__and4_1
XFILLER_21_175 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7517_ _7517_/D _7959_/RN _7958_/CLK _7517_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_147_350 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4729_ hold41/Z _4731_/A2 _4729_/B _7448_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_7448_ _7448_/D input75/Z _7589_/CLK _7448_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_174_37 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_135_567 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7379_ _7379_/D _7901_/RN _7810_/CLK _7379_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_116_770 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_107_20 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_130_250 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_89_698 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_88_175 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_67_24 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_130_272 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_29_231 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_57_551 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_177_2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_123_63 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_29_286 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_84_392 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_44_256 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_44_267 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_157_103 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_8_124 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_166_670 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_157_169 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_8_179 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_148_82 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_126_534 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_181_673 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_153_375 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_113_217 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_79_131 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_4_396 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_94_101 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_121_283 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_82_318 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_82_329 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_35_212 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_48_595 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_90_340 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_75_392 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_6750_ _7751_/Q _6644_/Z _6884_/B1 _7687_/Q _6752_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_63_587 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_63_576 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5701_ _5405_/B _5701_/A2 _5780_/A2 _5382_/Z _5701_/C _5702_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai221_2
XFILLER_92_2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3962_ input31/Z _4249_/A2 hold26/I _3961_/Z _3998_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_3893_ _7667_/Q _6039_/A1 _6022_/A1 _7659_/Q _6056_/A1 _7675_/Q _3896_/A1 VDD VSS
+ gf180mcu_fd_sc_mcu7t5v0__aoi222_2
X_6681_ _6681_/A1 _6681_/A2 _6681_/A3 _6681_/A4 _6684_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand4_1
XFILLER_148_147 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5632_ _5632_/A1 _5632_/A2 _5697_/A2 _5697_/A3 _5633_/A4 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor4_1
XFILLER_31_495 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5563_ _5663_/A1 _5405_/B _5381_/Z _5618_/B1 _5563_/B2 _5565_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai32_1
XFILLER_164_629 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_117_534 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7302_ input75/Z _4334_/Z _7302_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__and2_1
X_4514_ hold551/Z _4521_/A2 hold552/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
Xhold102 hold102/I _7416_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
XFILLER_172_673 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xhold135 hold135/I _7816_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
X_5494_ _5648_/A1 _5658_/B _5176_/B _5425_/B _5767_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_117_567 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xhold113 hold113/I hold113/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
Xhold124 hold124/I hold124/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
X_7233_ _7520_/Q _7233_/A2 _7233_/B1 _7518_/Q _7238_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_2
Xhold168 hold168/I hold168/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
Xhold146 hold146/I hold146/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
Xhold157 hold157/I _7565_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
X_4445_ hold761/Z _4487_/A1 _4450_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_4376_ _7214_/A1 _7214_/A2 _4376_/B _7511_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
Xhold179 hold179/I _6458_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
X_7164_ _7403_/Q _7203_/A2 _7204_/B1 _7389_/Q _7166_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_112_250 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6115_ hold73/Z _6123_/A2 _6115_/B _7695_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_86_602 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_451 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_440 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_98_495 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7095_ _7095_/A1 _7095_/A2 _7096_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_85_134 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_484 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_462 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_473 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_6046_ hold292/Z _6055_/A2 hold293/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_495 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2307 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2329 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2318 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1606 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_66_392 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_27_757 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_27_779 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7997_ _7997_/I _7997_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_1639 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1628 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1617 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_41_215 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_6948_ _6955_/A4 _6948_/A2 _6946_/Z _6948_/A4 _6949_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand4_4
XFILLER_179_283 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_10_602 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6879_ _6879_/A1 _6879_/A2 _6889_/C VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_10_613 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_167_478 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_148_670 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_108_534 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_163_651 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_150_334 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_104_740 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xhold680 _7472_/Q hold680/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
XFILLER_150_389 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xhold691 _7807_/Q hold691/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
XFILLER_131_570 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_77_602 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_1_377 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_89_495 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_94_33 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_92_605 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_92_627 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_64_318 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_17_212 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_94_88 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_91_137 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_33_716 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_13_451 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_43_92 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_43_81 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_43_70 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_145_139 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_9_499 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_154_662 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
Xoutput207 _3704_/ZN mgmt_gpio_oeb[8] VDD VSS gf180mcu_fd_sc_mcu7t5v0__buf_8
Xoutput218 _7992_/Z mgmt_gpio_out[18] VDD VSS gf180mcu_fd_sc_mcu7t5v0__buf_8
Xoutput229 _8002_/Z mgmt_gpio_out[28] VDD VSS gf180mcu_fd_sc_mcu7t5v0__buf_8
XFILLER_99_215 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_4230_ _7546_/Q _5807_/A1 _5871_/A1 _7582_/Q _4280_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_68_613 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_68_602 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_4_64 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4161_ _7669_/Q _6056_/A1 _4764_/A1 _7471_/Q _4162_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_122_592 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4092_ _4084_/Z _4092_/A2 _4092_/A3 _4092_/A4 _4107_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand4_2
XFILLER_83_627 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_82_126 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_67_189 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_7920_ _7920_/D _7961_/RN _7940_/CLK _7920_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
X_7851_ _7851_/D _7901_/RN _7851_/CLK _7851_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_48_392 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_6802_ _7433_/Q _7925_/Q _6802_/B1 _6802_/B2 _6804_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_4994_ _5602_/A2 _4993_/B _5648_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_2
X_7782_ _7782_/D _7901_/RN _7887_/CLK _7782_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffsnq_1
XFILLER_23_215 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_3945_ input50/Z _4275_/A2 _4231_/B1 input69/Z _3948_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_6733_ _7133_/S _6733_/A2 _6733_/B _7923_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_23_18 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_139_18 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6664_ _6878_/A2 _6664_/A2 _6664_/A3 _6880_/B1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor3_4
XFILLER_139_29 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5615_ _5689_/A1 _5692_/B _5618_/A3 _5763_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor3_1
X_3876_ _3796_/Z _4153_/A1 _5971_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_4
XFILLER_31_292 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_136_139 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6595_ _6599_/A2 _6618_/A3 _6596_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_5546_ _5797_/A2 _5546_/A2 _5546_/B1 _5543_/B _5546_/C _5646_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai221_2
X_5477_ _5496_/A1 _5797_/B _4965_/B _5543_/B _5477_/B2 _5510_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai32_1
XFILLER_2_108 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_7216_ _7216_/A1 _7216_/A2 _7941_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_4428_ _4428_/I _7963_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_160_676 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xclkbuf_2_3__f_mgmt_gpio_in[4] clkbuf_0_mgmt_gpio_in[4]/Z _4415_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_132_389 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_132_378 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_113_570 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7147_ _7683_/Q _7191_/A2 _6938_/I _7861_/Q _7148_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_59_635 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4359_ _4361_/A3 _4359_/A2 _4359_/B _7434_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_48_37 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_171_49 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7078_ _7210_/A2 _7078_/A2 _7078_/A3 _7078_/A4 _7078_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__or4_1
XFILLER_74_605 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_59_657 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6029_ hold181/Z _6038_/A2 hold182/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_46_318 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_58_189 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2115 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2126 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2104 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2159 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2148 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2137 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_104_98 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_1414 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1403 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_14_204 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_15_705 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1447 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1436 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1425 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_120_64 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1469 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1458 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_168_743 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_182_223 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_182_234 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_182_212 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_167_297 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_167_286 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_155_437 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_129_51 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_13_73 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_6_414 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_136_662 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_129_73 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_108_353 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_182_278 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_163_470 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_136_673 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_135_150 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_129_95 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_150_120 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_135_183 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_150_164 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_123_378 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_111_518 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_111_507 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_96_207 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_1_141 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_2_664 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_77_443 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_65_638 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_18_510 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_92_457 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_18_576 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_73_682 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_60_321 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_45_384 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1970 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_21_708 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1992 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1981 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_60_398 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_14_782 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_3730_ _7346_/Q _7345_/Q _3730_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_9_241 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3661_ _3661_/I _4368_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_173_212 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_159_798 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6380_ hold259/Z _6383_/A2 _6381_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_5400_ _5585_/A1 _5658_/B _5685_/B _5759_/A1 _5401_/A4 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_161_418 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5331_ _5645_/A1 _5687_/B _5618_/A3 _5331_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__or3_1
XFILLER_55_2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_141_131 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_142_676 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_5262_ _5687_/B _5504_/A3 _5779_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_114_367 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_7001_ _7605_/Q _6949_/I _7001_/B1 _7001_/B2 _7001_/C _7003_/B1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai221_1
X_5193_ _5199_/B _4915_/Z _4996_/Z _5202_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_114_389 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4213_ _7652_/Q _6022_/A1 _4843_/A1 _7507_/Q _4262_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_4144_ input44/Z _4275_/A2 hold108/I input62/Z _4198_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_56_605 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_95_273 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_18_29 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_28_318 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4075_ hold124/I _3963_/Z _4075_/B _4083_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_64_671 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7903_ _7903_/D _7961_/RN _7940_/CLK _7903_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
X_7834_ _7834_/D _7901_/RN _7834_/CLK _7834_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_63_170 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_51_321 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_7765_ _7765_/D _7901_/RN _7805_/CLK _7765_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_51_354 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4977_ _5603_/A1 _4993_/B _5669_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_4
X_6716_ _6716_/A1 _6716_/A2 _6716_/A3 _6716_/A4 _6721_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand4_1
X_3666__1 _3666__1/I _7279_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_3928_ _7796_/Q _6316_/A1 _3943_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_7696_ _7696_/D _7961_/RN _7704_/CLK _7696_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_20_741 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_149_286 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_109_106 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_3859_ hold146/Z hold118/Z _6158_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_4
X_6647_ _6878_/A2 _6665_/A2 _6665_/A3 _6647_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__and3_2
XFILLER_109_139 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6578_ _4352_/B _7907_/Q _6581_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_5529_ _5201_/B _5529_/A2 _5529_/A3 _5548_/A3 _5541_/A4 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand4_2
XFILLER_118_673 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_173_790 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_133_643 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_133_621 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_132_120 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_117_194 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_3_428 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_132_164 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_105_378 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_182_37 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_120_337 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_59_69 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_87_774 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_74_424 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_47_638 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_74_457 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_46_148 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_131_41 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_27_340 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_91_12 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1222 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1211 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1200 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_70_630 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_42_310 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_42_321 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_55_693 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_91_34 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1266 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1255 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1244 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1233 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_15_579 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1299 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1288 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1277 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_376 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_42_387 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_155_201 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_155_212 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_11_785 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_11_763 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_7_712 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_109_651 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_108_150 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_6_277 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_156_60 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_108_183 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_124_676 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_123_186 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_27_6 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_38_605 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_37_148 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_93_799 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_80_416 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_1_98 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_46_660 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4900_ _3722_/I _5006_/B _5006_/C _4900_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__and3_2
X_5880_ _4448_/Z _5880_/A2 _5880_/B _7585_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_92_298 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_61_641 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4831_ _4831_/A1 _7285_/A2 _4835_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_33_354 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_21_505 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_159_540 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_4762_ hold595/Z _4763_/A2 _4763_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_7550_ _7550_/D _7309_/Z _4418_/I1 _7550_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffnrnq_1
XFILLER_33_398 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_146_212 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4693_ hold161/Z _3819_/Z _4693_/B hold162/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_6501_ hold475/Z _6502_/A2 _6502_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_3713_ _7610_/Q _6826_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_7481_ _7481_/D _7944_/CLK _7481_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_6432_ hold68/Z _6434_/A2 _6432_/B _7844_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_3644_ _7411_/Q _4292_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__inv_3
XFILLER_161_215 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_134_418 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6363_ hold240/Z _6366_/A2 _6364_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_127_492 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_170_771 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6294_ hold47/Z _6298_/A2 _6294_/B _7779_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_130_602 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5314_ _5692_/B _5365_/B1 _5618_/A3 _5316_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor3_1
X_5245_ _3728_/I _5369_/B _5271_/A3 _5724_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor3_4
XFILLER_115_698 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
Xhold28 hold28/I hold28/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
Xhold17 hold17/I hold17/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
XFILLER_102_348 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xhold39 hold39/I hold39/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
X_5176_ _5027_/Z _5479_/A2 _5176_/B _5177_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_152_29 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_69_785 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_29_605 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_29_638 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_110_392 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_84_744 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4127_ _7749_/Q _6226_/A1 _4158_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_84_788 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_4058_ _4058_/A1 _4058_/A2 _4058_/A3 _4058_/A4 _4069_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor4_2
XFILLER_83_276 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_25_811 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_316 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_305 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_101_22 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_24_321 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7817_ _7817_/D _7901_/RN _7820_/CLK _7817_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XPHY_349 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_338 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_327 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_101_66 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_52_685 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_7748_ _7748_/D _7901_/RN _7810_/CLK _7748_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffsnq_1
XFILLER_137_212 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7679_ _7679_/D _7961_/RN _7704_/CLK _7679_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_165_543 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_152_259 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_106_676 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_105_120 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_133_495 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_86_12 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_126_85 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_120_134 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_86_34 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_120_156 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_47_402 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_101_392 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_74_232 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_28_660 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_90_747 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_90_736 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1030 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_43_641 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_96_9 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_70_471 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_70_460 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1074 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1063 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1052 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1041 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_140 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_43_674 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1096 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1085 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_156_510 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_168_392 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_129_779 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_167_70 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_167_81 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
Xhold509 _7860_/Q hold509/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
XFILLER_143_248 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_143_215 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_7_586 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_171_579 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_112_602 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_803 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_814 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_825 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_151_292 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5030_ _5496_/A1 _5458_/C _5661_/A1 _5031_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor3_1
XFILLER_111_123 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_97_357 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_836 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_847 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_858 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_869 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_18_2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_81_703 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_65_243 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6981_ _7709_/Q _7189_/A2 _7189_/B1 _7685_/Q _7189_/C1 _7653_/Q _6992_/A1 VDD VSS
+ gf180mcu_fd_sc_mcu7t5v0__aoi222_1
X_5932_ hold47/Z _5936_/A2 _5932_/B _7609_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_19_682 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_53_438 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_178_112 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5863_ hold355/Z _5868_/A2 _5864_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_21_302 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_167_808 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_7602_ _7602_/D _7901_/RN _7603_/CLK hold85/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
X_5794_ _5794_/A1 _5794_/A2 _5794_/A3 _5795_/A4 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand3_1
X_4814_ _4448_/Z _4816_/A2 _4814_/B _7494_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_166_318 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4745_ hold542/Z _4753_/S _4746_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_119_212 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_21_357 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7533_ _7533_/D _7961_/RN _7648_/CLK _7533_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_31_29 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4676_ _7463_/Q hold55/I hold48/Z hold49/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_7464_ _7464_/D _7901_/RN _7816_/CLK _7464_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_135_716 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6415_ hold68/Z _6417_/A2 _6415_/B _7836_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_7395_ _7395_/D _7961_/RN _7531_/CLK _7395_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
X_6346_ hold440/Z _6349_/A2 _6347_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
Xinput118 wb_adr_i[30] _4367_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
Xinput107 wb_adr_i[20] _5195_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_8
X_6277_ hold47/Z _6281_/A2 _6277_/B _7771_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
Xinput129 wb_dat_i[10] _7249_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_5228_ _5200_/B _3727_/I _3728_/I _5022_/B _5645_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand4_4
XFILLER_57_700 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5159_ _4965_/B _5366_/A2 _5797_/A2 _5752_/C VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor3_2
XFILLER_84_530 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_69_582 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_29_413 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_29_446 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_56_37 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_57_722 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_72_747 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_72_736 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_25_641 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_124 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_102 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_113 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_157 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_146 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_135 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_179 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_168 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_122_2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_180_321 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_125_237 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_125_215 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_4_534 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_21_73 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_180_354 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_137_73 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_4_589 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_121_432 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_79_357 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_87_390 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_47_210 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_48_744 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_47_232 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_90_566 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_71_780 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_4 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_176_605 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_16_696 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_148_318 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_30_176 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_30_187 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_129_576 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_129_565 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4530_ hold615/Z _4531_/A2 _4531_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_4461_ hold29/I hold6/Z hold7/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
Xhold317 _7379_/Q hold317/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
Xhold306 hold306/I _7795_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
XFILLER_7_97 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xclkbuf_leaf_100_csclk _7558_/CLK _7391_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_171_365 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_171_354 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xhold328 _7743_/Q hold328/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
XFILLER_116_259 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6200_ hold73/Z _6208_/A2 _6200_/B _7735_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
Xhold339 hold339/I _7659_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
X_7180_ _7960_/Q _7207_/A2 _7207_/B1 _7529_/Q _7205_/A2 _7533_/Q _7182_/A2 VDD VSS
+ gf180mcu_fd_sc_mcu7t5v0__aoi222_1
XFILLER_171_376 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6131_ hold423/Z _6140_/A2 _6132_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_600 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_4392_ _4392_/A1 _4396_/S _4393_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_97_121 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_611 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_622 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_633 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_100_605 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6062_ _4460_/Z _6072_/A2 _6062_/B hold208/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
XTAP_644 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_655 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_666 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_677 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_5013_ _5195_/B _4926_/Z _5010_/Z _5016_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor3_2
XTAP_688 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_699 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_26_29 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_38_276 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_54_736 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_54_747 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6964_ _7878_/Q _7203_/B1 _7193_/C1 _7724_/Q _6965_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_19_490 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_179_432 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5915_ hold47/Z hold276/Z _5915_/B _7601_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_34_460 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6895_ _6895_/A1 _6895_/A2 _6895_/A3 _6895_/A4 _6895_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__and4_1
X_5846_ _5846_/A1 _7285_/A2 _5848_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_166_104 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_21_132 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_166_137 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_5777_ _5777_/A1 _5777_/A2 _5777_/B _5777_/C _5802_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi211_2
X_7516_ _7516_/D _7959_/RN _7958_/CLK _7516_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
X_4728_ hold390/Z _4731_/A2 _4729_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_162_321 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4659_ hold55/I _4454_/Z hold36/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_108_738 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_107_226 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_107_215 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7447_ _7447_/D input75/Z _7447_/CLK _7447_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_162_354 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_135_557 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_7378_ _7378_/D _7901_/RN _7755_/CLK _7378_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
X_6329_ hold286/Z _6332_/A2 hold287/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_103_421 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_1_548 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_131_785 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_130_262 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_88_187 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_83_35 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_57_574 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_29_298 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_44_246 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_72_566 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_158_605 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xclkbuf_leaf_94_csclk _7558_/CLK _7573_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_53_780 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_12_132 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_40_463 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_13_688 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_12_187 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_12_176 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_148_72 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_181_641 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_153_354 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_114_719 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
Xclkbuf_leaf_32_csclk _7825_/CLK _7797_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
Xclkbuf_leaf_47_csclk clkbuf_3_7__f_csclk/Z _7821_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_94_157 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_48_530 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_94_179 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_36_747 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3961_ _7930_/Q _7578_/Q _7580_/Q _3961_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_16_460 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5700_ _5104_/B _5212_/Z _5780_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_149_627 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_149_638 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_148_115 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_3892_ _3892_/A1 _3892_/A2 _3892_/A3 _3892_/A4 _3918_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand4_2
X_6680_ _7716_/Q _6881_/A2 _6885_/A2 _7660_/Q _6681_/A4 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_5631_ _5331_/Z _5437_/B _5619_/Z _5697_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_85_2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_176_468 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5562_ _5735_/A2 _5585_/A1 _5562_/B _5704_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_163_129 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_157_682 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_144_321 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_129_373 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4513_ hold73/Z _4521_/A2 _4513_/B hold550/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_7301_ input75/Z _4334_/Z _7301_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__and2_1
X_7232_ _3658_/I _7281_/B1 _7233_/B1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
Xhold125 hold125/I _7750_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
X_5493_ _5603_/A1 _4993_/B _5797_/A2 _5493_/B _5530_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai31_1
Xhold114 hold114/I hold114/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
Xhold103 _7577_/Q hold103/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
Xhold136 _7808_/Q hold136/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
Xhold147 hold147/I _7718_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
Xhold158 _7706_/Q hold158/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
X_4444_ _4444_/A1 _7285_/A2 _4487_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_4
X_4375_ _4375_/A1 _4375_/A2 _7214_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_144_398 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
Xhold169 hold169/I _7439_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
X_7163_ _7407_/Q _7202_/A2 _7202_/B1 _7397_/Q _7385_/Q _7202_/C2 _7166_/A1 VDD VSS
+ gf180mcu_fd_sc_mcu7t5v0__aoi222_1
X_6114_ hold420/Z _6123_/A2 _6115_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_100_402 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_98_463 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_7094_ _7899_/Q _7197_/A2 _6938_/I _7859_/Q _7095_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XTAP_441 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_430 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_6045_ _4460_/Z _6055_/A2 _6045_/B hold254/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
XTAP_485 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_463 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_474 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_452 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_496 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2308 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_160_29 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2319 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_27_747 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_54_544 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_7996_ _7996_/I _7996_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_1629 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1618 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1607 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_169_16 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6947_ _7195_/A2 _7195_/C1 _7207_/B1 _7196_/B1 _6948_/A4 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor4_4
XFILLER_22_441 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_6878_ _7534_/Q _6878_/A2 _6879_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_50_761 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_167_424 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_139_126 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5829_ hold716/Z _5840_/A2 _5830_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_22_463 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_163_641 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_135_354 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_135_376 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_118_86 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
Xhold670 _7470_/Q hold670/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
XFILLER_1_312 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
Xhold681 _7531_/Q hold681/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
Xhold692 _7572_/Q hold692/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
XFILLER_134_41 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_103_295 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_94_67 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_76_179 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_18_747 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_72_374 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_60_558 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_9_423 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_9_412 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_41_783 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_139_682 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_126_321 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xoutput208 _3703_/ZN mgmt_gpio_oeb[9] VDD VSS gf180mcu_fd_sc_mcu7t5v0__buf_8
Xoutput219 _7993_/Z mgmt_gpio_out[19] VDD VSS gf180mcu_fd_sc_mcu7t5v0__buf_8
XFILLER_175_70 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_153_140 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_126_376 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_153_195 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_153_184 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_141_357 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_141_379 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4160_ _7653_/Q _6022_/A1 _4444_/A1 _7348_/Q _4779_/A1 _7477_/Q _4162_/A2 VDD VSS
+ gf180mcu_fd_sc_mcu7t5v0__aoi222_2
XFILLER_122_582 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_110_733 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_110_755 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4091_ _7638_/Q _5988_/A1 _4091_/B _4092_/A4 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_95_499 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_82_105 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7850_ _7850_/D _7901_/RN _7852_/CLK _7850_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
X_6801_ _7107_/A1 _6767_/C _7433_/Q _6802_/B2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_63_352 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_24_728 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7781_ _7781_/D _7901_/RN _7853_/CLK _7781_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
X_4993_ _5741_/A1 _5603_/A1 _4993_/B _4993_/C _4998_/C VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi211_1
X_3944_ _7892_/Q _6520_/A1 _4488_/A1 _7361_/Q _6209_/A1 _7746_/Q _3948_/A1 VDD VSS
+ gf180mcu_fd_sc_mcu7t5v0__aoi222_2
X_6732_ _7923_/Q _7133_/S _6733_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_3875_ _3886_/A2 hold133/Z _6384_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_4
X_6663_ _7910_/Q _7909_/Q _7908_/Q _6663_/A4 _6893_/C1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor4_4
X_5614_ _5614_/A1 _5642_/A2 _5614_/A3 _5614_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__and3_1
XFILLER_177_799 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6594_ _6586_/B _6594_/A2 _7910_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_5545_ _5662_/A1 _5545_/A2 _5545_/B _5764_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi21_2
XFILLER_145_641 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5476_ _5527_/A1 _5498_/A2 _5476_/B _5523_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_145_696 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_145_685 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_117_354 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7215_ _4376_/B _7511_/Q _7941_/Q _7215_/C _7216_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai211_1
X_4427_ _7413_/Q _4427_/A2 _4427_/B _4428_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_7146_ _7837_/Q _7203_/A2 _7193_/B1 _7635_/Q _7148_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_59_603 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_99_783 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_4358_ _7432_/Q _7581_/Q _4359_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_48_49 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_58_124 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_7077_ _7077_/A1 _7077_/A2 _7077_/A3 _7077_/A4 _7078_/A4 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand4_1
X_4289_ _7344_/Q _3734_/Z _7344_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_6028_ _4460_/Z _6038_/A2 _6028_/B hold201/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_86_499 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_58_179 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2105 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2116 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_104_88 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_73_149 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_54_330 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2149 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2138 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2127 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1415 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1404 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_70_812 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_64_37 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_1448 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1437 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1426 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_7979_ _7979_/D _7332_/Z _4418_/I1 _7979_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_2
XFILLER_54_396 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1459 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_558 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_167_232 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_80_25 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_10_411 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_23_783 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_168_788 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_155_405 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_22_271 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_129_41 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_129_63 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_108_321 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_135_195 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_97_709 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_151_688 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_123_357 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_2_676 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_150_176 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_150_187 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_145_73 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_49_157 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_161_50 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_77_499 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_64_105 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_18_500 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_61_812 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_33_503 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_45_352 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_45_363 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_72_171 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_33_514 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1960 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1993 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1982 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1971 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_159_777 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3660_ _3660_/I _4370_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_174_747 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_9_286 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_173_246 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_139_490 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_127_641 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_127_630 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_154_460 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5330_ _5200_/B _3727_/I _5369_/B _5648_/B2 _5335_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand4_1
XFILLER_181_290 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5261_ _5200_/B _3727_/I _5338_/A1 _5369_/B _5504_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand4_4
XFILLER_126_195 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_142_688 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_7000_ _6949_/I _6997_/Z _7000_/A3 _7000_/A4 _7001_/B2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand4_1
XFILLER_48_2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4212_ hold275/Z _4212_/A2 _5849_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_5192_ _5200_/B _5230_/A1 _5663_/A1 _5371_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor3_1
X_4143_ _4153_/A1 hold20/Z _4831_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_2
X_4074_ hold20/Z hold25/Z _5874_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_2
XFILLER_83_425 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_55_105 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_7902_ _7902_/D _7961_/RN _7940_/CLK _7902_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_70_108 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_36_352 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_48_190 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_52_812 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7833_ _7833_/D _7901_/RN _7883_/CLK _7833_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
X_7764_ _7764_/D _7901_/RN _7853_/CLK _7764_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_24_569 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_34_29 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4976_ _4993_/B _5604_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_6715_ _7760_/Q _6892_/A2 _6893_/C1 _7630_/Q _6716_/A4 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_51_388 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7695_ _7695_/D _7961_/RN _7735_/CLK _7695_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
X_3927_ _7940_/Q _7579_/Q _7580_/Q _3927_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_137_438 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3858_ hold146/Z hold113/Z _6282_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_4
X_6646_ _7910_/Q _6662_/A3 _6661_/A3 _6885_/B1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor3_4
X_3789_ _7337_/Q _7336_/Q _7414_/Q _3789_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_6577_ _7434_/Q _6590_/A1 _6586_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_173_780 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5528_ _3727_/I _5528_/A2 _5552_/A4 _5540_/B2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor3_2
XFILLER_152_408 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_133_611 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_145_493 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_160_463 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_160_452 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5459_ _5752_/B1 _5668_/A2 _5459_/B _5668_/B _5460_/A4 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XFILLER_132_132 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_105_357 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_59_48 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_132_176 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_120_316 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_99_580 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_7129_ _7129_/A1 _7129_/A2 _7129_/A3 _7128_/Z _7130_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand4_1
XFILLER_101_530 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_87_753 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_86_241 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_101_596 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_59_499 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_131_31 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_27_352 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_43_812 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1223 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1212 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1201 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_54_160 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_152_2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1256 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1245 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1234 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1289 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1278 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1267 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_156_747 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_156_725 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_11_753 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_6_201 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_156_758 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_155_246 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_109_641 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_171_739 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_7_779 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_6_256 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_108_195 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_151_496 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_111_305 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_78_742 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_172_60 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_93_723 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_93_712 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_65_425 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_65_436 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_93_778 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_18_374 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_34_812 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_45_160 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_52_108 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_178_316 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4830_ _7230_/A1 _4828_/S _4830_/B _7503_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
XTAP_1790 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_4761_ _4448_/Z _4763_/A2 _4761_/B _7468_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_4692_ _3819_/Z _4454_/Z _4693_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_3712_ _7609_/Q _7107_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_6500_ hold68/Z _6502_/A2 _6500_/B _7876_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_7480_ _7480_/D _7944_/CLK _7480_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_147_769 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3643_ _3643_/I _3801_/I0 VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_6431_ hold467/Z _6434_/A2 _6432_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_174_599 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_162_739 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_162_717 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6362_ hold47/Z _6366_/A2 _6362_/B _7811_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_161_238 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_155_780 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5313_ _5687_/C _5495_/B2 _5741_/B _5316_/C VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_170_761 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_142_463 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6293_ hold479/Z _6298_/A2 _6294_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_115_655 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_114_176 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5244_ _5779_/A1 _5433_/C _5273_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_69_720 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xhold29 hold29/I hold29/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
Xhold18 hold18/I hold18/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
X_5175_ _5749_/A2 _5175_/A2 _5178_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_84_701 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_28_105 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4126_ hold113/Z _3869_/I _4594_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_2
XFILLER_83_211 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4057_ _4057_/A1 _4057_/A2 _4057_/A3 _4057_/A4 _4058_/A4 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand4_1
XFILLER_71_428 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7816_ _7816_/D _7901_/RN _7816_/CLK _7816_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffsnq_1
XPHY_306 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_339 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_328 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_317 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_24_388 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_51_141 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7747_ _7747_/D _7901_/RN _7812_/CLK _7747_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
X_4959_ _5797_/B _4965_/B _5774_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_4
XFILLER_101_89 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_7678_ _7678_/D _7901_/RN _7819_/CLK _7678_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffsnq_1
XFILLER_138_747 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6629_ _6634_/A1 _7906_/Q _6659_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_153_728 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_118_460 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_3_215 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_133_441 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_161_783 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_121_647 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_120_179 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_75_712 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_19_73 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_47_425 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_75_778 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_16_812 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_34_108 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_1031 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1020 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_15_344 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1064 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1053 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1042 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1097 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1086 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1075 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_175_319 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_30_358 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_128_213 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_156_588 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_109_460 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_137_780 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_124_463 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_804 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_815 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_826 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_837 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_848 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_859 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_25_4 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_93_531 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_93_575 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6980_ _7376_/Q _7188_/A2 _6990_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_5931_ hold413/Z _5936_/A2 _5932_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_53_428 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_81_759 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_80_247 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_179_636 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5862_ _4460_/Z _5868_/A2 _5862_/B _7577_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_33_152 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_33_141 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7601_ _7601_/D _7901_/RN _7821_/CLK hold57/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
X_5793_ _5104_/B _5793_/A2 _5793_/B _5794_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_61_494 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4813_ hold682/Z _4816_/A2 _4814_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_178_179 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4744_ _4448_/Z _4753_/S _4744_/B _7458_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_7532_ _7532_/D _7961_/RN _7532_/CLK _7532_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
X_7463_ _7463_/D _7901_/RN _7463_/CLK _7463_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
X_4675_ hold55/I hold47/Z hold48/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_135_706 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6414_ hold508/Z _6417_/A2 _6415_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_7394_ _7394_/D input75/Z _7573_/CLK _7394_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_162_558 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6345_ hold47/Z _6349_/A2 _6345_/B _7803_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_143_783 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6276_ hold484/Z _6281_/A2 _6277_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_103_603 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xinput108 wb_adr_i[21] _5302_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_4
XFILLER_170_591 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_142_282 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5227_ _5199_/B _5201_/B _5338_/A1 _5369_/B _5573_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor4_4
XFILLER_102_124 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
Xinput119 wb_adr_i[31] _4367_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_102_179 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_88_369 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_69_572 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_57_712 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5158_ _5496_/A1 _5527_/A1 _5167_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_2
XFILLER_29_425 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_29_436 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5089_ _3728_/I _5022_/B _5303_/A3 _5285_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_84_542 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4109_ _4206_/A1 _7223_/A1 _4109_/B _4110_/I0 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_57_789 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_16_108 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_112_99 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_72_37 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_125 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_24_141 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_25_686 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_103 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_114 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_169_146 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_158 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_147 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_136 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_25_697 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_169_168 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_169 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_12_347 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_8_318 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_8_329 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_181_812 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_119_780 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_115_2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_180_344 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_153_558 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_141_709 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_134_761 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_106_463 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_97_56 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_106_496 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_94_317 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_752 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_153_73 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_153_84 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_121_499 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_121_488 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_75_586 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_35_428 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_90_534 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_62_247 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_71_770 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_15_141 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_5 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_16_686 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_87_6 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_31_678 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_169_691 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_172_812 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_7_32 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4460_ hold29/Z hold6/Z _4460_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__and2_4
Xhold307 _7711_/Q hold307/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
XFILLER_144_525 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_7_373 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
Xhold329 _7728_/Q hold329/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
Xhold318 _7632_/Q hold318/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
X_4391_ _4387_/S _7889_/Q _4391_/B _4391_/ZN VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_2
XFILLER_125_783 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6130_ _4460_/Z _6140_/A2 _6130_/B hold211/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_140_753 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_140_742 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_140_731 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_124_271 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_601 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_612 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_623 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_634 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_30_2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_97_144 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_6061_ hold207/Z _6072_/A2 _6062_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_58_509 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_645 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_656 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_667 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_5012_ _4926_/Z _5010_/Z _5195_/B _5139_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_4
XFILLER_85_339 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_678 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_689 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_38_200 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_38_211 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_39_712 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_66_531 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_66_586 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6963_ _7870_/Q _7195_/C1 _7207_/B1 _7716_/Q _6965_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_179_422 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5914_ hold57/Z hold276/I _5915_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_81_567 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_22_601 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6894_ _7400_/Q _6894_/A2 _6659_/Z _7471_/Q _6894_/C1 _7404_/Q _6895_/A4 VDD VSS
+ gf180mcu_fd_sc_mcu7t5v0__aoi222_1
XFILLER_53_269 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5845_ _4454_/Z _5845_/A2 _5845_/B _7570_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_179_499 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_179_488 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_21_144 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_42_29 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_166_127 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_158_29 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5776_ _5776_/A1 _5778_/A1 _5776_/A3 _5776_/A4 _5777_/C VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand4_1
XFILLER_163_812 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7515_ _7515_/D _7959_/RN _7958_/CLK _7515_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_108_717 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4727_ hold73/Z _4731_/A2 _4727_/B _7447_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_4658_ _7425_/Q _4685_/A1 _4661_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_147_374 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_107_205 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_7446_ _7446_/D input75/Z _7589_/CLK _8006_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_123_709 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xinput90 spimemio_flash_io2_oeb input90/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_7377_ _7377_/D _7901_/RN _7755_/CLK _7377_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffsnq_1
XFILLER_116_761 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_88_100 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4589_ _4589_/A1 _7285_/A2 _4593_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_6328_ hold47/Z _6332_/A2 _6328_/B hold306/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_131_764 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_6259_ hold468/Z _6264_/A2 _6260_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_103_499 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_76_317 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_67_59 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_123_32 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_17_428 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_123_98 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_72_534 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_72_589 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_25_450 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_13_645 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_40_442 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_9_638 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_172_108 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_154_812 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_32_51 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_32_73 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_166_683 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_126_525 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_4_321 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_107_783 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_121_241 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_79_144 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_82_309 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_593 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3960_ hold630/I hold107/Z hold108/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_4
XFILLER_51_729 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_73_80 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_149_617 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_148_105 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3891_ _7619_/Q _5937_/A1 _4488_/A1 _7362_/Q _3892_/A4 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_43_280 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5630_ _5776_/A1 _5778_/A1 _5697_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_148_149 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5561_ _5741_/A1 _4993_/B _5663_/A1 _5561_/B _5562_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai31_1
XFILLER_78_2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_156_160 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_145_812 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5492_ _5648_/A1 _5735_/A2 _5685_/B _5648_/B2 _5642_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_129_363 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_8_671 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4512_ hold548/Z _4521_/A2 hold549/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_7300_ input75/Z _4334_/Z _7300_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__and2_1
X_7231_ _7281_/A2 _3658_/I _7233_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_171_130 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xhold115 hold115/I _7377_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
Xhold104 _7539_/Q hold104/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
Xhold126 _7540_/Q hold126/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
XFILLER_171_141 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4443_ hold11/Z hold31/Z _7506_/Q hold32/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_4
Xhold137 _7792_/Q hold137/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
XFILLER_104_219 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
Xhold148 _7606_/Q hold148/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
Xhold159 hold159/I _6138_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
X_4374_ _4906_/S _4374_/A2 _4374_/A3 _4374_/A4 _4375_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand4_1
X_7162_ _7525_/Q _7190_/C1 _7168_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_6113_ _4460_/Z _6123_/A2 _6113_/B hold203/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_7093_ _7891_/Q _7196_/A2 _7196_/B1 _7641_/Q _7095_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_86_615 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_442 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_431 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_420 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_6044_ hold253/Z _6055_/A2 _6045_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_86_637 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_464 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_475 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_453 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_100_447 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_100_436 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_497 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_486 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_85_169 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_73_309 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2309 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_7995_ _7995_/I _7995_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_54_534 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1619 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1608 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_6946_ _6946_/A1 _6946_/A2 _6946_/A3 _6946_/A4 _6946_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__and4_1
XFILLER_26_247 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_41_239 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_22_431 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6877_ _7133_/S _6877_/A2 _6877_/B _7929_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_167_436 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_139_116 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5828_ _5828_/A1 _7285_/A2 _5840_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_4
X_5759_ _5759_/A1 _5768_/A3 _5779_/A2 _5779_/A1 _5759_/C _5760_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi221_1
XFILLER_154_108 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_147_171 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_136_812 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_147_193 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_135_333 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7429_ hold50/Z _7901_/RN _7450_/CLK _7986_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_135_366 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_2_803 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_162_196 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xhold660 _7383_/Q hold660/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
Xhold671 _7570_/Q hold671/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
XFILLER_1_302 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xhold693 _7629_/Q hold693/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
Xhold682 _7494_/Q hold682/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
XFILLER_1_357 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_76_125 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_94_24 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_182_2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_94_57 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_18_715 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_72_331 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_27_73 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_45_567 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_60_548 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_40_250 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_127_801 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_173_417 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_173_428 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xclkbuf_3_7__f_csclk clkbuf_0_csclk/Z clkbuf_3_7__f_csclk/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_127_812 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_5_641 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_181_461 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_114_528 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_114_517 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_99_206 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xoutput209 _4405_/Z mgmt_gpio_out[0] VDD VSS gf180mcu_fd_sc_mcu7t5v0__buf_8
XFILLER_126_388 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_5_696 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_4_44 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_4090_ _4090_/A1 _4090_/A2 _4090_/A3 _4091_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_64_810 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_82_139 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_36_534 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6800_ _6800_/A1 _6800_/A2 _6800_/A3 _6799_/Z _6802_/B1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand4_1
XFILLER_91_651 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_36_556 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4992_ _5254_/A2 _5608_/A1 _4993_/C VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_4
X_7780_ _7780_/D _7901_/RN _7797_/CLK _7780_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_23_206 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_51_515 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_177_712 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_3943_ _3943_/A1 _3943_/A2 _3943_/A3 _3943_/A4 _3954_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand4_2
X_6731_ _7433_/Q _7922_/Q _6731_/B1 _6731_/B2 _6733_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_176_211 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_149_425 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3874_ _3835_/Z hold133/Z _6333_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_4
X_6662_ _7910_/Q _6663_/A4 _6662_/A3 _6892_/B1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor3_4
X_5613_ _5359_/B _5613_/A2 _5678_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_149_469 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_31_283 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_164_417 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_136_108 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_118_812 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6593_ _7434_/Q _6767_/C _6593_/B1 _7910_/Q _6594_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_5544_ _5547_/A1 _5547_/A2 _5651_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_129_193 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5475_ _5066_/Z _5680_/A1 _5475_/B _5502_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_7214_ _7214_/A1 _7214_/A2 _7517_/D _7216_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_4426_ _7412_/Q _7415_/Q _4427_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_7145_ _7829_/Q _7202_/A2 _7205_/B1 _7747_/Q _7148_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_98_250 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_101_712 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4357_ _7433_/Q _4361_/A2 _4359_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
Xclkbuf_leaf_93_csclk _7558_/CLK _7871_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_58_103 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_171_29 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7076_ _7818_/Q _7207_/A2 _7207_/B1 _7720_/Q _7076_/C _7077_/A4 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi221_1
XFILLER_86_456 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4288_ _7345_/Q _4288_/A2 _7345_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XFILLER_104_34 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_104_23 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_101_778 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6027_ hold200/Z _6038_/A2 _6028_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_73_117 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2106 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2117 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_67_692 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_27_534 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2139 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2128 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1405 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_82_673 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_27_567 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_27_556 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1438 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1427 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1416 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_81_150 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_14_206 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_42_515 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7978_ _7978_/D _7331_/Z _4418_/I1 _7978_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_54_375 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_54_386 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_154_6 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
Xclkbuf_leaf_31_csclk clkbuf_3_7__f_csclk/Z _7806_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_120_44 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_120_33 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1449 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_6929_ _6953_/A1 _6950_/A1 _6941_/A2 _7189_/C1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor3_4
XFILLER_80_37 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_22_250 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_23_795 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_155_428 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_109_812 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_182_247 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xclkbuf_leaf_46_csclk clkbuf_3_7__f_csclk/Z _7583_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_89_13 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_170_409 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_135_163 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_135_141 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_129_86 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_163_494 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_123_314 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_8_2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_150_133 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
Xhold490 hold490/I _4472_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
XFILLER_89_283 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_150_199 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_161_73 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_18_534 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_159_712 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1961 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1950 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_72_183 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_158_211 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1994 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1983 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1972 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_60_389 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_41_570 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_13_283 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_9_221 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_118_108 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_9_298 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5260_ _5199_/B _5201_/B _3728_/I _5022_/B _5768_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor4_4
XFILLER_114_325 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_142_656 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_141_144 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4211_ hold146/I _4075_/B _5855_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_5191_ _5476_/B _5689_/A2 _5191_/B1 _5191_/B2 _7520_/Q _5362_/B1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai221_1
XFILLER_110_531 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4142_ _7677_/Q _6073_/A1 _4174_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_68_434 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_110_564 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4073_ _4427_/B _4073_/A2 _4073_/A3 _4073_/B _7551_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai31_1
XFILLER_95_286 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7901_ _7901_/D _7901_/RN _7901_/CLK _7901_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_83_459 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_64_651 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_7832_ _7832_/D _7901_/RN _7883_/CLK _7832_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffsnq_1
XFILLER_64_673 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_63_150 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_24_526 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4975_ _5069_/A2 _4930_/Z _4953_/Z _4975_/A4 _4993_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand4_4
X_7763_ _7763_/D _7901_/RN _7805_/CLK _7763_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_91_492 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_149_200 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_6714_ _7816_/Q _6880_/A2 _6891_/B1 _7670_/Q _6716_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_3926_ hold25/Z _4155_/A2 hold26/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_4
X_7694_ _7694_/D _7961_/RN _7694_/CLK _7694_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffsnq_1
XFILLER_137_428 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3857_ _4075_/B _4217_/A2 _4444_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_4
X_6645_ _7910_/Q _6664_/A3 _6658_/A3 _6882_/B1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor3_4
XFILLER_50_29 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_166_29 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_164_247 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_149_299 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3788_ _3801_/S hold144/Z hold52/Z _3925_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi21_4
XFILLER_118_620 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_20_798 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_6576_ _6634_/A1 _6633_/A2 _6658_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_4
X_5527_ _5527_/A1 _5689_/A2 _5548_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_117_141 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_172_291 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5458_ _5496_/A1 _5527_/A1 _5458_/B _5458_/C _5668_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi211_2
XFILLER_132_122 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_117_196 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_105_347 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_99_570 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5389_ _5705_/A2 _5585_/A1 _5624_/B _5759_/A1 _5736_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_4409_ input1/Z _7607_/Q _4409_/B _4409_/ZN VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_2
X_7128_ _6949_/I _7128_/A2 _7128_/A3 _7128_/A4 _7128_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__and4_1
XFILLER_115_88 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_115_77 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7059_ _7680_/Q _7191_/A2 _7190_/B1 _7616_/Q _7190_/A2 _7794_/Q _7063_/A1 VDD VSS
+ gf180mcu_fd_sc_mcu7t5v0__aoi222_1
XFILLER_74_404 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_39_191 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_131_65 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_131_54 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1213 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1202 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_312 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1257 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1246 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1235 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1224 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_70_632 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_54_183 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_145_2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1279 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1268 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_70_676 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_42_389 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_168_531 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_23_570 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_156_737 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_7_703 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_151_453 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_123_144 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_2_463 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_27_8 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_172_83 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_78_798 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_92_201 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_77_286 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_77_275 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_92_256 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_73_470 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_65_70 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_45_150 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_46_673 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_178_328 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1780 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1791 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_14_581 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_4760_ hold679/Z _4763_/A2 _4761_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_119_428 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4691_ _7437_/Q _4718_/A1 _4694_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_3711_ _7608_/Q _7079_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_174_534 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_146_247 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3642_ hold51/I _5640_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_6430_ hold47/Z _6434_/A2 _6430_/B _7843_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_6361_ hold268/Z _6366_/A2 _6362_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_60_2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5312_ _5724_/B _5624_/A2 _5741_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_170_751 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6292_ hold41/Z _6298_/A2 _6292_/B _7778_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_5243_ _5714_/B1 _5687_/B _5247_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_2
Xhold19 hold19/I hold19/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
X_5174_ _5735_/A2 _5643_/A2 _5027_/Z _5643_/B1 _5175_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_69_776 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_69_765 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_29_607 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4125_ hold113/Z _3881_/Z _4554_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_2
XFILLER_83_223 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_56_437 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_4056_ _7623_/Q _5954_/A1 _5988_/A1 _7639_/Q _4057_/A4 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_45_29 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XPHY_307 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_101_13 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7815_ _7815_/D _7961_/RN _7815_/CLK _7815_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffsnq_1
XFILLER_24_334 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_52_643 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_329 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_318 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_12_507 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_52_676 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4958_ _4941_/C _4941_/B _4973_/A3 _4920_/Z _4965_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai22_4
X_7746_ _7746_/D _7901_/RN _7746_/CLK _7746_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
X_3909_ _7354_/Q _4444_/A1 _6124_/A1 _7707_/Q _3911_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_7677_ _7677_/D _7961_/RN _7702_/CLK _7677_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffsnq_1
XFILLER_20_540 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_20_551 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4889_ hold674/Z _4892_/A2 _4890_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_6628_ _7921_/Q _7133_/S _6686_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_165_567 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_4_717 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_106_623 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6559_ _7902_/Q _6559_/A2 _6560_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_105_144 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_160_250 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_126_32 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_10_65 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_121_637 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_87_540 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_87_551 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_86_69 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_47_404 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_59_286 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_19_106 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_142_53 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_90_749 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_90_727 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_28_673 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1021 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_27_183 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_1010 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1065 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1054 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1032 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1043 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_35_73 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_1098 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1087 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1076 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_128_203 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_156_534 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_128_247 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_7_566 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_112_615 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_111_103 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_805 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_816 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_151_283 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_3_783 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_827 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_838 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_849 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_66_735 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_65_212 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_81_716 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5930_ hold41/Z _5936_/A2 _5930_/B _7608_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_7600_ _7600_/D _7901_/RN _7673_/CLK _7600_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_80_259 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5861_ hold103/Z _5868_/A2 _5862_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_34_676 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5792_ _7545_/Q _5520_/C _5792_/B1 _5792_/B2 _5806_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_4812_ _4812_/A1 _7285_/A2 _4816_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_166_309 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4743_ hold76/Z _4753_/S _4744_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_7531_ _7531_/D _7961_/RN _7531_/CLK _7531_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
X_7462_ _7462_/D _7901_/RN _7463_/CLK _7462_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
X_4674_ _7986_/I _4685_/A1 _4677_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_147_567 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_135_718 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_107_409 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6413_ hold47/Z _6417_/A2 _6413_/B _7835_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_7393_ _7393_/D input75/Z _7573_/CLK _7393_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_134_239 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_6344_ hold419/Z _6349_/A2 _6345_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_115_442 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_143_795 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_142_250 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6275_ hold41/Z _6281_/A2 _6275_/B _7770_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
Xinput109 wb_adr_i[22] _5224_/A4 VDD VSS gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_170_581 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5226_ _5006_/C _5616_/A1 _5433_/C _5290_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_130_456 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_111_692 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5157_ _5179_/B _5783_/A2 _5173_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_57_724 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5088_ _5338_/A1 _5369_/B _5054_/Z _5114_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor3_4
XFILLER_96_392 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_84_565 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_84_554 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4108_ _7549_/Q _4206_/A1 _4109_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_29_448 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_57_779 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_84_598 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_84_576 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_71_215 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_4039_ _4039_/I0 _7552_/Q _4427_/B _7552_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_24_120 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_72_49 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_24_131 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_40_602 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_104 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_115 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_148 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_137 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_126 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_52_495 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_7729_ _7729_/D _7901_/RN _7753_/CLK _7729_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_166_810 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_157_309 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_159 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_12_337 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_178_692 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_138_534 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_20_392 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_165_386 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_4_514 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_4_525 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_153_548 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_125_239 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_108_2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_180_389 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_161_570 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_137_86 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_97_46 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_79_304 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_133_283 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_121_434 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_47_212 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_101_191 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_63_705 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_47_223 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_75_565 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_6 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_16_676 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_30_101 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_175_139 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_129_567 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xhold308 _7627_/Q hold308/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
Xhold319 hold319/I _7632_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
X_4390_ _4387_/S input90/Z _4391_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_124_250 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_98_602 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_140_721 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_602 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_613 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_624 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_635 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_646 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_657 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_668 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_6060_ _4454_/Z _6072_/A2 _6060_/B _7669_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_5011_ _5211_/A3 _5011_/A2 _5011_/B _5016_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi21_2
XFILLER_66_510 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_23_2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_679 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_78_392 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_66_576 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_38_256 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_6962_ _7894_/Q _7197_/A2 _7189_/C1 _7652_/Q _6965_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_53_215 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_179_412 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5913_ hold41/Z hold276/Z _5913_/B _7600_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_6893_ _7402_/Q _6893_/A2 _6893_/B1 _7390_/Q _6893_/C1 _7473_/Q _6895_/A3 VDD VSS
+ gf180mcu_fd_sc_mcu7t5v0__aoi222_1
X_5844_ hold671/Z _5845_/A2 _5845_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_61_292 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_166_117 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7514_ _7514_/D _7959_/RN _7958_/CLK _7514_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
X_5775_ _5775_/A1 _5775_/A2 _5801_/A1 _5786_/C1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_147_331 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_147_342 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_4726_ hold494/Z _4731_/A2 _4727_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_174_172 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4657_ _4685_/A1 hold77/Z _4657_/B hold78/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_135_515 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_107_217 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7445_ _7445_/D input75/Z _7447_/CLK _7445_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_174_29 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_7376_ _7376_/D _7901_/RN _7746_/CLK _7376_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffsnq_1
Xinput91 spimemio_flash_io3_do input91/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
Xinput80 spi_sck input80/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_162_389 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6327_ hold304/Z _6332_/A2 hold305/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_107_12 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_101_9 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4588_ _4454_/Z _4588_/A2 _4588_/B _7398_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_143_570 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_131_721 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_115_283 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6258_ hold41/Z _6264_/A2 _6258_/B _7762_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_5209_ _5209_/A1 _5209_/A2 _5209_/A3 _5376_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand3_2
X_6189_ hold68/Z _6191_/A2 _6189_/B _7730_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_88_189 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_29_212 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_123_44 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_123_77 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_123_88 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_60_719 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_16_64 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_25_495 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_52_270 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_8_105 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_166_662 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_40_498 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_148_74 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_5_801 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_32_85 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_4_333 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_106_250 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_107_795 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_164_95 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_121_231 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_121_286 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_95_638 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_90_321 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_75_384 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_35_215 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_44_760 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_73_70 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3890_ _7382_/Q hold114/I _6452_/A1 _7861_/Q _3892_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_176_459 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5560_ _5613_/A2 _5560_/A2 _5590_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_129_353 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5491_ _5542_/A2 _5542_/A3 _5517_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_157_684 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4511_ _4460_/Z _4521_/A2 _4511_/B hold233/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_4442_ hold11/Z _3810_/S _4442_/B hold12/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi21_4
Xhold105 _3792_/Z _3795_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
Xhold116 _7544_/Q hold116/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
X_7230_ _7230_/A1 _7228_/S _7230_/B _7949_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_7_160 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_172_676 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
Xhold138 hold138/I _6322_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
Xhold127 _3790_/Z hold127/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
Xhold149 hold149/I _5926_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
X_4373_ _4925_/A1 _4923_/A1 _4365_/Z _4374_/A4 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor3_1
XFILLER_144_389 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_125_570 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7161_ _7133_/S _7161_/A2 _7161_/A3 _7161_/B _7938_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai31_1
X_6112_ hold202/Z _6123_/A2 _6113_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_98_454 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_86_605 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7092_ _7649_/Q _7195_/A2 _7195_/B1 _7625_/Q _7195_/C1 _7875_/Q _7097_/A3 VDD VSS
+ gf180mcu_fd_sc_mcu7t5v0__aoi222_1
XTAP_432 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_421 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_410 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_6043_ _4454_/Z _6055_/A2 _6043_/B hold586/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_140_595 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_86_627 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_58_318 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_465 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_476 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_454 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_443 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_112_297 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_100_459 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_498 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_487 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_7994_ _7994_/I _7994_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_1609 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_81_354 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6945_ _7189_/C1 _7190_/B1 _7196_/A2 _7193_/C1 _6946_/A4 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor4_1
XFILLER_169_18 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6876_ _7929_/Q _7133_/S _6877_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_50_752 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_179_275 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_179_286 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_10_605 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_5827_ hold41/Z _5827_/A2 _5827_/B _7562_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_5758_ _5614_/Z _5758_/A2 _5758_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_148_662 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_4709_ hold57/Z _3819_/Z _4709_/B hold58/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_147_183 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_118_33 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5689_ _5689_/A1 _5689_/A2 _5757_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_7428_ hold44/Z _7901_/RN _7450_/CLK _7985_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_162_153 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_135_378 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_118_44 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_162_186 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
Xhold650 _7748_/Q hold650/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
XFILLER_89_421 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_89_410 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_78_37 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_7359_ _7359_/D _7961_/RN _7875_/CLK _7359_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
Xhold661 _7399_/Q hold661/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
Xhold672 _7524_/Q hold672/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
Xhold694 _7847_/Q hold694/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
Xhold683 _7509_/Q hold683/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
XFILLER_134_32 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_131_562 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_89_487 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_89_476 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_77_638 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_134_87 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_103_286 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_92_619 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_175_2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_72_321 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_17_215 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_57_373 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_33_708 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_60_516 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_26_782 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_13_421 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_9_425 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_9_414 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_43_73 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_159_73 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_9_469 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_126_334 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_154_676 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_153_186 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_107_570 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_4_34 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_122_540 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_68_605 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_67_126 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_391 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_95_479 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_83_608 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_48_384 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_91_641 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_63_354 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4991_ _5206_/A2 _5136_/A1 _5585_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_4
X_6730_ _7027_/A1 _6767_/C _7433_/Q _6731_/B2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_3942_ _7353_/Q _4444_/A1 _4249_/A2 input32/Z _3943_/A4 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_2
XFILLER_90_2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3873_ _3796_/Z hold118/Z _6107_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_4
X_6661_ _6878_/A2 _6662_/A3 _6661_/A3 _6894_/C1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor3_4
X_5612_ _5599_/Z _5612_/A2 _5610_/Z _5639_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand3_1
X_6592_ _6618_/A3 _6830_/B _6593_/B1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_164_407 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5543_ _5741_/A3 _5545_/A2 _5543_/B _5543_/C _5547_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XFILLER_8_480 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_160_602 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_145_687 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_144_131 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_144_142 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_5474_ _5461_/Z _5474_/A2 _5474_/B _5521_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_7213_ _7133_/S _7213_/A2 _7213_/B _7940_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_4425_ _7979_/Q _4425_/A2 _4425_/ZN VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_2
X_7144_ _7140_/Z _7144_/A2 _7144_/A3 _7144_/A4 _7159_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand4_1
X_4356_ _6937_/A1 _6953_/A1 _6950_/A1 _4361_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor3_1
XFILLER_113_584 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_99_774 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_86_402 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_48_29 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_140_392 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_7075_ _7075_/A1 _7075_/A2 _7075_/A3 _7076_/C VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_101_757 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4287_ _7346_/Q _4287_/A2 _7346_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XFILLER_74_619 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6026_ _4454_/Z _6038_/A2 _6026_/B _7653_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
XTAP_2107 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_39_373 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_54_321 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2129 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2118 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1406 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_66_192 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1439 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1428 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1417 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_7977_ _7977_/D _7330_/Z _7977_/CLK _7977_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_42_527 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6928_ _7914_/Q _7913_/Q _6937_/A1 _6599_/Z _7200_/B1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor4_4
XFILLER_54_398 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_167_212 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_147_6 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_23_752 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6859_ _6859_/A1 _6859_/A2 _6859_/A3 _6860_/C VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_6_406 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_129_43 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_136_676 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_150_112 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_145_20 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_108_389 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_1_100 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xhold480 _7350_/Q hold480/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
XFILLER_2_656 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
Xhold491 hold491/I _7351_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
XFILLER_1_144 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_77_424 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_38_73 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_38_84 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_73_641 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_45_354 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_73_696 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_33_505 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_45_376 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_1951 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1940 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_54_61 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1995 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1984 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1973 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1962 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_60_379 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_41_560 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_173_215 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_173_248 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_182_760 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_142_602 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_127_698 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_126_175 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4210_ _7586_/Q _5881_/A1 _4754_/A1 _7466_/Q _4243_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_5190_ _5424_/A1 _5680_/B2 _5755_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_122_392 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4141_ hold118/Z hold107/Z _4873_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_68_457 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4072_ _7551_/Q _4427_/B _4073_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_95_90 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7900_ _7900_/D _7901_/RN _7900_/CLK _7900_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_36_321 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_36_354 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_48_181 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_91_482 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7831_ _7831_/D _7901_/RN _7887_/CLK _7831_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffsnq_1
X_4974_ _5201_/B _5210_/A3 _4974_/A3 _5797_/C VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand3_4
X_7762_ _7762_/D _7901_/RN _7868_/CLK _7762_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_177_521 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_149_212 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3925_ hold123/Z _3925_/A2 hold127/Z _3794_/Z _4155_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand4_4
X_6713_ _7702_/Q _6889_/A2 _6887_/B1 _7678_/Q _6659_/Z _7622_/Q _6716_/A2 VDD VSS
+ gf180mcu_fd_sc_mcu7t5v0__aoi222_1
X_7693_ _7693_/D _7961_/RN _7701_/CLK _7693_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffsnq_1
XFILLER_51_357 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_51_368 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_177_532 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_149_234 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_20_733 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_6644_ _7910_/Q _6665_/A2 _6659_/A3 _6644_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__and3_2
XFILLER_177_587 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_177_576 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3856_ hold19/Z _3787_/Z hold127/Z _3794_/Z _4217_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand4_4
X_3787_ hold51/Z hold144/Z _3801_/S _3787_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_4
X_6575_ _7907_/Q _7906_/Q _6590_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_2
XFILLER_180_708 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_164_259 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5526_ _5066_/Z _5680_/B2 _5552_/A4 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_118_676 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5457_ _5741_/A3 _5099_/B _5776_/A1 _3723_/I _5457_/C _5459_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai221_1
XFILLER_105_337 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_59_39 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4408_ input1/Z input2/Z _4409_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_182_29 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_120_318 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5388_ _5772_/A1 _5614_/A1 _5783_/C VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_4339_ _7518_/Q _4438_/A2 _7513_/Q _4340_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_7127_ _7754_/Q _7201_/A2 _7205_/B1 _7746_/Q _7128_/A4 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_101_532 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7058_ _7133_/S _7058_/A2 _7058_/A3 _7058_/B _7934_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai31_1
XFILLER_86_298 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6009_ _4454_/Z _6021_/A2 _6009_/B _7645_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_28_811 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_55_641 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_82_460 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1214 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1203 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_70_611 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_27_354 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_54_140 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_91_26 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_82_482 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_82_493 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_1247 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1236 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1225 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_168_521 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1269 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1258 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_11_700 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_42_368 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_138_2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_155_226 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_155_248 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_155_215 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_10_276 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_124_602 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_6_247 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_124_613 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_156_85 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_104_392 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_78_744 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_92_246 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_18_321 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_18_332 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_18_387 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_178_318 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1770 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_33_357 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1781 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1792 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_81_70 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_60_176 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xclkbuf_leaf_92_csclk _7558_/CLK _7587_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
X_3710_ _7623_/Q _3710_/ZN VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_159_565 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4690_ _4718_/A1 hold165/Z _4690_/B hold166/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_3641_ _7540_/Q _5522_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_6360_ hold41/Z _6366_/A2 _6360_/B _7810_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_5311_ _5645_/A1 _5687_/B _5624_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_4
XFILLER_115_602 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_53_2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6291_ hold501/Z _6298_/A2 _6292_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_115_657 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_130_605 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5242_ _5689_/A1 _5563_/B2 _5575_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_102_318 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5173_ _5476_/B _5498_/A2 _5173_/B _5173_/C _5178_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai211_1
Xclkbuf_leaf_30_csclk clkbuf_3_7__f_csclk/Z _7799_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_84_703 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_68_243 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4124_ hold20/Z hold133/Z _4579_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_84_747 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xinput1 debug_mode input1/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_56_427 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xclkbuf_leaf_45_csclk clkbuf_3_7__f_csclk/Z _7603_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
X_4055_ input38/Z _5903_/A1 _5971_/A1 _7631_/Q _4057_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_37_641 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_64_493 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_36_173 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_36_195 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_7814_ _7814_/D _7961_/RN _7815_/CLK _7814_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffsnq_1
XPHY_319 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_308 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_40_806 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_51_154 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_52_666 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4957_ _5069_/A2 _4930_/Z _4953_/Z _4957_/A4 _5797_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand4_4
X_7745_ _7745_/D _7901_/RN _7812_/CLK _7745_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_61_29 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_177_373 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_131_9 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_7676_ _7676_/D _7901_/RN _7821_/CLK _7676_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffsnq_1
X_3908_ _7747_/Q _6209_/A1 _4232_/A2 input10/Z _3911_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_4888_ _4888_/A1 _7285_/A2 _4892_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_137_215 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3839_ _3817_/I hold113/Z _6299_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_4
X_6627_ _6556_/B _7002_/B _7133_/S VDD VSS gf180mcu_fd_sc_mcu7t5v0__and2_4
XFILLER_137_248 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6558_ _7433_/Q _4331_/Z _6562_/A1 _4352_/B _6564_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_2
XFILLER_106_602 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5509_ _5509_/A1 _5509_/A2 _5505_/Z _5509_/A4 _5519_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor4_1
XFILLER_126_11 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_106_635 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6489_ hold708/Z _6502_/A2 _6490_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_120_126 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_86_37 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_87_596 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_59_276 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_75_758 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_83_780 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_15_302 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_16_803 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_83_791 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1022 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1000 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1011 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_70_463 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_1055 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1033 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1044 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_15_357 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_1099 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1088 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1077 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1066 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_176 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_129_705 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_156_546 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_171_505 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_167_73 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_51_73 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_112_605 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_2_250 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_806 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_817 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_124_498 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_111_115 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_828 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_839 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_120_671 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_120_660 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_78_596 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_66_747 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_19_641 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_38_449 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_46_460 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_53_408 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_5860_ hold73/Z _5868_/A2 _5860_/B _7576_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_18_195 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_179_638 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_73_290 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_22_806 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4811_ _7230_/A1 _4809_/S _4811_/B _7493_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
XTAP_2290 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_5791_ _5691_/Z _5791_/A2 _5760_/Z _5791_/A4 _5792_/B2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand4_1
XFILLER_61_496 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_61_474 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4742_ hold55/Z _4742_/A2 _4753_/S VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_4
X_7530_ _7530_/D _7961_/RN _7642_/CLK _7530_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
X_7461_ _7461_/D _7901_/RN _7461_/CLK _7461_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_174_321 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4673_ _4685_/A1 hold43/Z _4673_/B hold44/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_119_215 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_174_343 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_147_579 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6412_ hold523/Z _6417_/A2 _6413_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_128_771 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7392_ _7392_/D _7901_/RN _7887_/CLK _7392_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_115_410 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6343_ hold41/Z _6349_/A2 _6343_/B _7802_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_6274_ hold386/Z _6281_/A2 _6275_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_209 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5225_ _5563_/B2 _5687_/B _5624_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_4
XFILLER_103_638 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_102_104 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_130_446 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_69_552 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_5156_ _5600_/A1 _5797_/B _5797_/A2 _5542_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor3_1
XFILLER_130_479 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_111_682 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_56_29 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5087_ _4898_/Z _5777_/A1 _5087_/B _5087_/C _5094_/B1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai211_1
X_4107_ _4107_/A1 _4107_/A2 _4107_/A3 _7223_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor3_4
XFILLER_84_544 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_25_600 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4038_ _4284_/A1 _4807_/A1 _4038_/B _4039_/I0 VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_112_68 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_65_780 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_105 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_116 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_149 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_138 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_127 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_12_316 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5989_ hold746/Z _6004_/A2 _5990_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_24_187 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_24_176 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_52_463 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_7728_ _7728_/D _7901_/RN _7813_/CLK _7728_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_165_354 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7659_ _7659_/D _7961_/RN _7735_/CLK _7659_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_153_505 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_137_54 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xoutput190 _3685_/ZN mgmt_gpio_oeb[27] VDD VSS gf180mcu_fd_sc_mcu7t5v0__buf_8
XFILLER_0_776 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_47_202 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_153_97 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_102_693 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_48_747 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_7 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_55_290 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_94_9 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_71_783 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_31_636 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_156_321 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_62_83 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_30_179 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_11_382 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_171_302 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_144_538 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_7_89 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
Xhold309 hold309/I _7627_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
XFILLER_171_357 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_140_744 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_3_570 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_603 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_614 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_625 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_5010_ _5200_/B _5201_/B _5230_/A1 _5024_/A2 _5010_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__or4_4
XTAP_636 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_647 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_658 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_97_168 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_669 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_38_202 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_78_382 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_66_544 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_16_2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6961_ _7822_/Q _7202_/A2 _7196_/B1 _7636_/Q _7196_/A2 _7886_/Q _6967_/A2 VDD VSS
+ gf180mcu_fd_sc_mcu7t5v0__aoi222_1
XFILLER_47_780 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5912_ hold172/Z hold276/I _5913_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_6892_ _7386_/Q _6892_/A2 _6892_/B1 _7532_/Q _6895_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_5843_ _4448_/Z _5845_/A2 _5843_/B _7569_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_34_463 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_167_619 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_10_809 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_21_124 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_7513_ _7513_/D _7959_/RN _7958_/CLK _7513_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
X_5774_ _5774_/A1 _5774_/A2 _5774_/B1 _5774_/B2 _5774_/C _5801_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi221_2
XFILLER_175_641 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_159_192 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_147_354 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4725_ _4460_/Z _4731_/A2 _4725_/B hold109/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_4656_ hold76/Z hold55/Z _4656_/B hold77/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_7444_ _7444_/D input75/Z _7447_/CLK _7444_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
X_7375_ _7375_/D _7901_/RN _7852_/CLK _7375_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffsnq_1
Xinput70 mgmt_gpio_in[7] input70/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
Xinput81 spi_sdo input81/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_4587_ hold613/Z _4588_/A2 _4588_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_6326_ hold41/Z _6332_/A2 _6326_/B _7794_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_116_763 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xinput92 spimemio_flash_io3_oeb input92/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_89_603 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_107_24 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_89_647 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6257_ hold499/Z _6264_/A2 _6258_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_115_295 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_107_68 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_107_79 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_67_28 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5208_ _5015_/B _5197_/Z _5392_/A2 _5709_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor3_2
X_6188_ hold252/Z _6191_/A2 _6189_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_88_179 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_5139_ _5139_/A1 _5014_/Z _5209_/A1 _5498_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand3_2
XFILLER_97_691 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_72_503 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_53_783 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_13_647 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_12_124 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_138_321 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_12_179 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_165_140 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_120_2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_153_357 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_180_176 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_122_733 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_4_389 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_122_744 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_122_788 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_94_105 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_562 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_57_50 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_91_812 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_75_352 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_48_566 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_90_344 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_51_709 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_16_463 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_157_641 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_129_332 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_31_488 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_31_499 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_172_611 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_172_600 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5490_ _5543_/B _5498_/A2 _5497_/A3 _5542_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor3_1
XFILLER_156_140 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_8_673 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_8_662 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4510_ hold231/Z _4521_/A2 hold232/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_4441_ hold31/I _7506_/Q _4442_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__and2_1
Xhold117 _3805_/Z hold117/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
Xhold139 hold139/I _7792_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
X_7160_ _7611_/Q _7210_/A2 _7160_/B _7433_/Q _7161_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi211_1
Xhold128 _3847_/Z hold128/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
X_4372_ _4372_/A1 _4372_/A2 _4372_/A3 _4372_/A4 _4375_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand4_1
X_6111_ _4454_/Z _6123_/A2 _6111_/B _7693_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
XTAP_400 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_7091_ _7697_/Q _7194_/A2 _7194_/B1 _7665_/Q _7194_/C1 _7811_/Q _7097_/A2 VDD VSS
+ gf180mcu_fd_sc_mcu7t5v0__aoi222_1
XTAP_433 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_422 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_411 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_6042_ hold584/Z _6055_/A2 hold585/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_112_254 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_86_617 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_455 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_466 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_444 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_499 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_488 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_477 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_82_812 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_54_503 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7993_ _7993_/I _7993_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_94_694 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_93_171 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_66_385 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6944_ _7195_/B1 _7194_/B1 _7203_/B1 _7200_/B1 _6946_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor4_1
XFILLER_54_558 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_35_783 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6875_ _7433_/Q _7928_/Q _6875_/B1 _6875_/B2 _6877_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_5826_ hold483/Z _5827_/A2 _5827_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_5757_ _5425_/B _5757_/A2 _5757_/B _5783_/B _5758_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XFILLER_182_419 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_182_408 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_175_460 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_163_611 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_4708_ _3819_/Z hold47/Z _4709_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_162_121 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5688_ _5705_/B _5555_/B _5688_/A3 _5725_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor3_1
XFILLER_108_549 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7427_ hold75/Z _7901_/RN _7450_/CLK _7984_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
X_4639_ hold63/Z _3830_/Z _4639_/B hold64/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_135_357 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_162_176 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xhold662 _8002_/I hold662/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
Xhold640 _7855_/Q hold640/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
X_7917__346 _7917_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__tieh
Xhold651 _7476_/Q hold651/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
X_7358_ _7358_/D _7961_/RN _7587_/CLK _7358_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffsnq_2
Xhold673 _7660_/Q hold673/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
XFILLER_104_744 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6309_ hold41/Z _6315_/A2 _6309_/B _7786_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
Xhold695 _7564_/Q hold695/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
X_7289_ _4454_/Z _7289_/A2 _7289_/B _7961_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
Xhold684 _7546_/Q hold684/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
XFILLER_103_276 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_89_499 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_76_105 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_94_37 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_85_694 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_168_2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_27_64 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_150_98 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_158_449 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_139_641 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_13_499 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_40_263 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_166_471 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_166_460 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_138_140 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_175_51 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_181_496 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_175_73 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_153_176 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_122_530 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_110_747 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_95_425 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_82_108 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_64_812 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_48_330 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_48_341 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_36_525 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4990_ _5394_/A1 _5254_/A2 _5136_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_2
XFILLER_90_174 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_17_783 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3941_ _7852_/Q _6435_/A1 _6265_/A1 _7772_/Q _3943_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_51_539 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_177_736 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3872_ _3886_/A2 hold118/Z _6124_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_4
X_6660_ _7910_/Q _6664_/A2 _6664_/A3 _6884_/B1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor3_4
X_5611_ _5672_/A2 _5606_/B _5749_/A4 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_83_2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6591_ _7910_/Q _6879_/A1 _6767_/C VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_4
X_5542_ _5166_/B _5542_/A2 _5542_/A3 _5542_/A4 _5542_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__or4_1
XFILLER_117_302 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_172_463 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5473_ _5473_/A1 _5473_/A2 _5776_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_117_357 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_144_187 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_144_176 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_117_379 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7212_ _7940_/Q _7133_/S _7213_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_4424_ _4424_/A1 input73/Z _4424_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__and2_1
X_7143_ _7813_/Q _7194_/C1 _7204_/A2 _7845_/Q _7144_/A4 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_99_753 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_4355_ _7912_/Q _6599_/A2 _6950_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_4
X_7074_ _7752_/Q _7201_/A2 _7201_/B1 _7672_/Q _7075_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_58_105 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4286_ _7345_/Q _7344_/Q _3734_/Z _4287_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_104_14 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_67_650 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6025_ hold718/Z _6038_/A2 _6026_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_2108 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_104_47 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_82_620 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_39_363 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_55_812 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2119 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_70_804 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_64_29 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_15_709 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_27_558 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_54_344 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_54_355 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_120_13 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1429 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1418 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1407 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_81_141 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_42_517 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7976_ _7976_/D _7329_/Z _4418_/I1 _7976_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
X_6927_ _6950_/A1 _6955_/A4 _6908_/Z _7194_/C1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor3_4
XFILLER_80_39 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_23_775 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6858_ _7494_/Q _6882_/B1 _6647_/Z _7468_/Q _6859_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_168_747 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_10_403 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_50_572 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5809_ _4448_/Z _5811_/A2 _5809_/B _7546_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_148_460 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6789_ _7665_/Q _6885_/A2 _6647_/Z _7617_/Q _6887_/B1 _7681_/Q _6791_/A2 VDD VSS
+ gf180mcu_fd_sc_mcu7t5v0__aoi222_1
XFILLER_136_666 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_129_88 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_163_496 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_2_602 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_150_146 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
Xhold470 _7861_/Q hold470/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
Xhold481 hold481/I _4467_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
XFILLER_2_646 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_150_179 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
Xhold492 _7664_/Q hold492/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
XFILLER_49_116 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_64_108 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_85_491 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_61_804 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_45_344 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_1952 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1941 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1930 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1985 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1974 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1963 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1996 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_9_212 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_158_257 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_167_780 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_70_83 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_126_143 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_182_772 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_154_463 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_126_187 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_141_146 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_79_70 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_68_414 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4140_ hold20/Z hold113/Z _4584_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_96_756 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_1_690 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_110_566 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_95_266 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4071_ _7550_/Q _4206_/A1 _4073_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_83_428 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_37_812 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7830_ _7830_/D _7901_/RN _7834_/CLK _7830_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffsnq_1
XFILLER_63_130 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_4973_ _3727_/I _4920_/Z _4973_/A3 _4975_/A4 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor3_2
X_7761_ _7761_/D _7901_/RN _7873_/CLK _7761_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
X_6712_ _7734_/Q _6878_/A2 _6712_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__or2_1
X_7692_ _7692_/D _7961_/RN _7692_/CLK _7692_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffsnq_1
X_3924_ input9/Z _4232_/A2 _3940_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_6643_ _7910_/Q _6663_/A4 _6664_/A2 _6881_/B1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor3_4
XFILLER_165_728 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3855_ _3817_/I hold133/Z _6435_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_4
X_3786_ _7506_/Q hold51/Z hold52/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__and2_1
X_6574_ _6633_/A2 _6618_/A3 _6574_/B _7906_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_5525_ _5543_/C _5498_/B _5545_/A2 _5542_/A4 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor3_1
XFILLER_117_132 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_173_783 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_160_411 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5456_ _5087_/B _5456_/A2 _5433_/C _5457_/C VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_105_327 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_121_809 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_59_29 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4407_ _7607_/Q _4334_/Z _4407_/B _4407_/ZN VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_2
X_5387_ _5600_/A1 _5797_/B _4993_/C _5618_/A3 _5409_/B2 _5587_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai32_1
XFILLER_132_179 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_87_712 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4338_ _5903_/A2 _4338_/A2 _4338_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__or2_1
X_7126_ _7820_/Q _7207_/A2 _7207_/B1 _7722_/Q _7205_/A2 _7738_/Q _7128_/A3 VDD VSS
+ gf180mcu_fd_sc_mcu7t5v0__aoi222_1
XFILLER_59_425 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_59_436 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_7057_ _7934_/Q _7133_/S _7058_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_4269_ _7862_/Q _6469_/A1 _6537_/A1 _7894_/Q _4271_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_28_801 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6008_ hold636/Z _6021_/A2 _6009_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_46_108 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_131_23 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1204 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_7959_ _7959_/D _7959_/RN _4411_/I1 hold31/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_131_89 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1248 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1237 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1226 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1215 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1259 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_70_667 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_24_32 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_145_4 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_11_712 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_155_205 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_7_716 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_24_87 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_149_780 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_11_778 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_7_727 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_171_709 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_109_655 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_151_411 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_136_463 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_124_669 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_151_455 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_123_168 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_151_499 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_78_734 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_49_73 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_77_277 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_65_428 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_19_812 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_73_450 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_61_601 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_45_141 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_46_664 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_60_100 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1760 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_21_509 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1782 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1793 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1771 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_3640_ _7539_/Q _5362_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_155_783 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_127_463 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6290_ hold73/Z _6298_/A2 _6290_/B _7777_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_5310_ _5687_/C _5495_/B2 _5550_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_154_282 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_127_496 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5241_ _5199_/B _5201_/B _4915_/Z _5433_/C _5623_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand4_2
XFILLER_114_146 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_69_712 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_46_2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5172_ _5669_/A1 _5027_/Z _5173_/C VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_114_179 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_96_531 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_69_767 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4123_ hold113/Z _4151_/A2 _4564_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_4054_ _7671_/Q _6056_/A1 _6209_/A1 _7743_/Q _4057_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_1
Xinput2 debug_oeb input2/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_28_108 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_83_225 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xclkbuf_opt_1_0_csclk _7961_/CLK clkbuf_opt_1_0_csclk/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
X_7813_ _7813_/D _7901_/RN _7813_/CLK _7813_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_101_15 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_24_336 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7744_ _7744_/D _7901_/RN _7746_/CLK _7744_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XPHY_309 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_101_37 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_101_26 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_51_144 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4956_ _4944_/Z _4956_/A2 _5602_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_2
XFILLER_52_689 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_177_363 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_7675_ _7675_/D _7961_/RN _7691_/CLK _7675_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
X_3907_ input28/Z _4239_/A2 hold134/I _7821_/Q _3911_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_20_531 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4887_ _4454_/Z _4887_/A2 _4887_/B _7534_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_3838_ _3850_/A1 _3864_/A2 _3843_/A3 hold274/I hold113/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand4_4
X_6626_ _7001_/C _7434_/Q _7002_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_2
XFILLER_153_709 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6557_ _6557_/I _6559_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_3769_ _7968_/Q _7969_/Q _3772_/S _7969_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_5508_ _5765_/A2 _5508_/A2 _5649_/A3 _5509_/A4 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_118_463 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_10_34 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6488_ _4448_/Z _6502_/A2 _6488_/B _7870_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_126_34 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5439_ _5727_/A2 _5439_/A2 _5439_/A3 _5439_/A4 _5445_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand4_1
XFILLER_105_168 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_133_499 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_133_488 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_120_105 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7109_ _7133_/S _7109_/A2 _7109_/B _7936_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_142_33 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_47_428 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_74_236 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_74_247 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_19_98 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_27_141 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_55_461 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_55_494 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1001 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1012 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_150_2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1056 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1034 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1045 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1023 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_70_475 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1089 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1078 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1067 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_30_317 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_171_517 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_137_783 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_7_579 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_136_282 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_109_496 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_3_763 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_807 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_111_127 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_3_785 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_818 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_829 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_120_650 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_93_567 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_81_718 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_81_707 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_74_770 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_46_450 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_19_697 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_179_628 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_178_105 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2280 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_33_144 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_34_656 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4810_ _7493_/Q _4809_/S _4811_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_2291 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_5790_ _5790_/A1 _5790_/A2 _5791_/A4 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_175_812 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4741_ hold559/Z _4753_/I1 _4741_/S _4741_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XTAP_1590 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_7460_ hold10/Z _7901_/RN _7461_/CLK hold9/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
X_4672_ _7462_/Q hold55/I hold42/Z hold43/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_147_536 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6411_ hold41/Z _6417_/A2 _6411_/B _7834_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_128_761 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7391_ _7391_/D _7901_/RN _7391_/CLK _7391_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_115_422 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6342_ hold388/Z _6349_/A2 _6343_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_115_444 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_88_306 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6273_ hold73/Z _6281_/A2 _6273_/B _7769_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_5224_ _5302_/A1 _5195_/B _5224_/A3 _5224_/A4 _5687_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__or4_4
XFILLER_142_263 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_115_499 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5155_ _5774_/A1 _5643_/A2 _5155_/B _5769_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_69_586 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_29_428 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_56_203 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5086_ _5648_/A1 _5087_/B _5682_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_4106_ _4106_/A1 _4106_/A2 _4106_/A3 _4106_/A4 _4107_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand4_2
XFILLER_84_534 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_56_247 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4037_ _7551_/Q _4284_/A1 _4038_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_112_58 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_71_239 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_37_494 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_72_29 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_13_807 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_24_122 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_106 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_52_431 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_139 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_128 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_117 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
X_5988_ _5988_/A1 _7285_/A2 _6004_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_4
XFILLER_40_615 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_4939_ _4900_/Z _4915_/Z _5199_/B _4973_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi21_4
X_7727_ _7727_/D _7901_/RN _7813_/CLK _7727_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_166_812 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7658_ _7658_/D _7961_/RN _7694_/CLK _7658_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_177_193 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6609_ _6953_/A1 _6609_/A2 _6611_/A2 _6908_/A1 _7914_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai22_1
XFILLER_165_366 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_119_783 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_119_761 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7589_ _7589_/D input75/Z _7589_/CLK _7999_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_21_33 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_180_336 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_137_44 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_134_731 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_4_538 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_161_561 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_97_37 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_121_425 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_106_477 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xoutput180 _3694_/ZN mgmt_gpio_oeb[18] VDD VSS gf180mcu_fd_sc_mcu7t5v0__buf_8
Xoutput191 _3684_/ZN mgmt_gpio_oeb[28] VDD VSS gf180mcu_fd_sc_mcu7t5v0__buf_8
XFILLER_0_733 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_744 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
Xclkbuf_leaf_91_csclk _7558_/CLK _7370_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_75_567 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_62_239 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_16_601 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_56_770 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_71_762 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_15_144 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XPHY_8 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_16_667 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_43_453 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_102_80 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_70_250 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_31_626 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_43_464 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_62_51 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_157_812 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_156_388 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_7_354 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_7_365 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
Xclkbuf_leaf_44_csclk clkbuf_3_7__f_csclk/Z _7450_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_152_550 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_98_615 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_98_626 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_98_637 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_3_560 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_604 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_615 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_112_458 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_87_70 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xclkbuf_leaf_59_csclk clkbuf_3_6__f_csclk/Z _7704_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XTAP_626 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_637 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_648 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_659 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_94_810 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_66_501 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_66_534 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_93_353 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6960_ _7692_/Q _7194_/A2 _7188_/A2 _7375_/Q _7782_/Q _7202_/B1 _6967_/A1 VDD VSS
+ gf180mcu_fd_sc_mcu7t5v0__aoi222_1
XFILLER_38_247 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5911_ hold73/Z hold276/Z _5911_/B _7599_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_47_792 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_62_751 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_19_494 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6891_ _7408_/Q _6891_/A2 _6891_/B1 _7508_/Q _6891_/C1 _7394_/Q _6895_/A1 VDD VSS
+ gf180mcu_fd_sc_mcu7t5v0__aoi222_1
X_5842_ hold764/Z _5845_/A2 _5843_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_5773_ _5658_/B _5606_/B _5773_/B _5773_/C _5775_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XFILLER_61_283 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7512_ _7512_/D _7959_/RN _7958_/CLK _7517_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_166_108 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_148_812 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4724_ _8006_/I _4731_/A2 _4725_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_147_333 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_147_366 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_4655_ hold55/Z _4448_/Z _4656_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_7443_ hold93/Z _7961_/RN _7603_/CLK _7443_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
Xinput60 mgmt_gpio_in[31] input60/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
Xinput71 mgmt_gpio_in[8] input71/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
Xinput82 spi_sdoenb _3663_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_7374_ _7374_/D _7961_/RN _7573_/CLK _7374_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
X_4586_ _4448_/Z _4588_/A2 _4586_/B _7397_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_143_550 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_6325_ hold315/Z _6332_/A2 _6326_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_116_753 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_116_742 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
Xinput93 trap input93/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_131_723 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_131_712 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_107_36 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_103_425 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6256_ hold73/Z _6264_/A2 _6256_/B _7761_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_103_458 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5207_ _5203_/I _5207_/A2 _5392_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_6187_ hold47/Z _6191_/A2 _6187_/B _7729_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_5138_ _4365_/Z _5138_/A2 _5209_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_111_491 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_96_191 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_57_567 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5069_ _4906_/Z _5069_/A2 _5210_/B _5069_/A4 _5458_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand4_4
XFILLER_84_375 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_45_729 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_80_570 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_52_250 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_139_812 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_178_491 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_32_43 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_181_634 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_119_591 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_119_580 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_113_2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_107_775 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_121_222 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_48_534 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_91_802 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_57_73 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_71_570 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_44_762 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_71_581 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_31_434 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_43_294 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_148_108 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_31_478 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
Xhold107 _3959_/Z hold107/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
X_4440_ input75/Z _4334_/Z _4440_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_171_144 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xhold129 hold129/I _7710_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
XFILLER_144_347 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
Xhold118 hold118/I hold118/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
X_4371_ _4922_/A3 _4922_/A4 _4924_/A1 _4924_/A2 _4374_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor4_1
XFILLER_171_177 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_125_572 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_113_712 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_113_701 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6110_ hold723/Z _6123_/A2 _6111_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_140_531 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7090_ _7851_/Q _7193_/A2 _7193_/B1 _7633_/Q _7193_/C1 _7729_/Q _7097_/A1 VDD VSS
+ gf180mcu_fd_sc_mcu7t5v0__aoi222_1
XTAP_423 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_401 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_412 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_6041_ _4448_/Z _6055_/A2 _6041_/B _7660_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_140_575 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_98_467 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_58_309 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_456 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_467 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_445 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_434 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_79_692 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_489 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_478 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_39_534 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_39_545 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_39_567 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7992_ _7992_/I _7992_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_94_673 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_81_312 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_26_206 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6943_ _7194_/A2 _7189_/B1 _7201_/B1 _7190_/C1 _6946_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor4_1
XFILLER_54_548 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_179_211 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_81_378 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_34_250 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6874_ _7184_/A1 _6767_/C _7433_/Q _6875_/B2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_5825_ hold73/Z _5827_/A2 _5825_/B _7561_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_167_428 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5756_ _5756_/A1 _5756_/A2 _5756_/A3 _7543_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__or3_1
XFILLER_147_141 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4707_ _7441_/Q _4718_/A1 _4710_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_5687_ _5689_/A1 _5689_/A2 _5687_/B _5687_/C _5688_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi211_1
X_4638_ _3830_/Z hold41/Z _4639_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_7426_ hold56/Z _7901_/RN _7450_/CLK _7983_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_163_667 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
Xhold630 hold630/I hold630/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
Xhold641 _7462_/Q hold641/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
XFILLER_162_166 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
Xhold652 _7740_/Q hold652/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
XFILLER_116_583 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
Xhold663 _7767_/Q hold663/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
X_7357_ _7357_/D _7961_/RN _7370_/CLK _7357_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffsnq_2
X_4569_ _4569_/A1 _7285_/A2 _4573_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
Xhold685 _7676_/Q hold685/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
XFILLER_104_756 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6308_ hold369/Z _6315_/A2 _6309_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_7288_ hold773/Z _7289_/A2 _7289_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
Xhold696 _7466_/Q hold696/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
Xhold674 _7535_/Q hold674/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
X_6239_ hold251/Z _6242_/A2 _6240_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_134_34 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_94_16 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_990 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_57_353 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_72_323 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_72_389 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_13_401 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_25_283 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_41_743 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_53_570 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_158_406 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_159_53 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_43_75 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_159_97 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_5_611 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_153_144 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_4_176 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_4_58 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_76_673 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3940_ _3940_/A1 _3940_/A2 _3940_/A3 _3940_/A4 _3954_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand4_2
XFILLER_63_378 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_16_250 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_32_743 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_44_570 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_149_428 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3871_ _4212_/A2 hold113/Z _6316_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_4
XFILLER_32_776 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_176_247 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5610_ _5602_/Z _5610_/A2 _5610_/A3 _5609_/Z _5610_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__and4_1
XFILLER_31_286 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6590_ _6590_/A1 _6665_/A2 _6879_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_2
XFILLER_176_269 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5541_ _5369_/B _5024_/Z _5543_/B _5541_/A4 _5550_/C VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor4_2
XFILLER_129_141 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_118_804 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_76_2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_145_634 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_129_163 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_8_460 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5472_ _5668_/A2 _5462_/Z _5472_/B _5472_/C _5474_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XFILLER_105_509 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_7211_ _7433_/Q _7939_/Q _7211_/B _7213_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_4423_ input85/Z input58/Z _7980_/Q _4423_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_7142_ _7789_/Q _7202_/B1 _7205_/A2 _7739_/Q _7144_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_4354_ _6908_/A1 _7913_/Q _6953_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_4
X_7073_ _7736_/Q _7205_/A2 _7205_/B1 _7744_/Q _7075_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_101_704 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_59_607 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_140_383 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4285_ _7344_/Q _3734_/Z _4288_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_6024_ _4448_/Z _6038_/A2 _6024_/B _7652_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_100_247 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_39_353 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_104_37 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_100_269 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_73_109 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2109 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_7975_ _7975_/D _7328_/Z _7977_/CLK _7975_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XTAP_1419 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1408 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_82_676 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_81_164 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6926_ _6937_/A1 _6951_/A2 _7203_/B1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_4
XFILLER_120_25 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_35_570 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6857_ _7527_/Q _6885_/B1 _6890_/A2 _7474_/Q _6859_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_50_540 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_167_247 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6788_ _7803_/Q _6883_/A2 _6883_/B1 _7787_/Q _6791_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_5808_ hold684/Z _5811_/A2 _5809_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_5739_ _5739_/A1 _5739_/A2 _5739_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_136_601 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_109_804 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_13_34 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_6_408 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_135_100 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_108_314 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_135_144 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7409_ _7409_/D _7901_/RN _7876_/CLK _7409_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_145_22 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xhold460 _7764_/Q hold460/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
Xhold471 _7773_/Q hold471/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
XFILLER_104_531 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_150_158 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_145_55 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
Xhold493 hold493/I _7664_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
XFILLER_77_404 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
Xhold482 hold482/I _7350_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
XFILLER_89_286 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_1_168 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_49_106 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_38_53 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_46_802 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_180_2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_58_673 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_58_695 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_18_526 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_72_120 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_72_142 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1942 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1931 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1920 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_73_698 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_72_175 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_60_337 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1986 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1975 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1964 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1953 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_13_242 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_158_247 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1997 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_14_798 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_13_286 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_167_792 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_167_770 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_139_483 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_139_494 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_182_795 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
Xclkbuf_2_2__f_mgmt_gpio_in[4] clkbuf_0_mgmt_gpio_in[4]/Z _4031_/C2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_181_283 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_5_496 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_5_485 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_110_534 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_95_212 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_68_426 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4070_ _4284_/A1 _7224_/I0 _4073_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_95_70 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_64_676 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_7760_ _7760_/D _7901_/RN _7868_/CLK _7760_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffsnq_1
X_4972_ _5006_/C _5608_/A1 _5714_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_2
XFILLER_17_570 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_36_389 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3923_ _7828_/Q _6384_/A1 _6418_/A1 _7844_/Q _3943_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_7691_ _7691_/D _7961_/RN _7691_/CLK _7691_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
X_6711_ _7686_/Q _6884_/B1 _6716_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_3854_ hold124/Z hold113/Z _6226_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_4
X_6642_ _6878_/A2 _7909_/Q _7908_/Q _6663_/A4 _6882_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor4_4
XFILLER_32_573 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_177_589 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_177_567 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3785_ hold143/Z _7337_/Q _7414_/Q _3785_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_9_780 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6573_ _7434_/Q _6633_/A2 _6574_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_5524_ _5524_/I _5558_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_118_667 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_117_144 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_172_250 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_160_401 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_145_486 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_132_103 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5455_ _5648_/A2 _4996_/Z _5643_/A2 _5705_/A2 _5657_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_133_637 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4406_ _7963_/Q _4334_/Z _4407_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_7125_ _7780_/Q _7200_/A2 _7201_/B1 _7674_/Q _7200_/B1 _7868_/Q _7128_/A2 VDD VSS
+ gf180mcu_fd_sc_mcu7t5v0__aoi222_1
X_5386_ _5669_/B _5669_/A1 _5292_/B _5621_/B _5716_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_4337_ _5903_/A2 _4338_/A2 _4438_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_115_25 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_99_584 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_115_69 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_113_394 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_101_567 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_87_768 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_86_256 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_86_245 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7056_ _7001_/C _7933_/Q _7058_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_4268_ _7692_/Q _6107_/A1 _4769_/A1 _7472_/Q _4271_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_75_29 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_6007_ _4448_/Z _6021_/A2 _6007_/B _7644_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_4199_ _7887_/Q _6520_/A1 _5988_/A1 _7637_/Q _5841_/A1 _7570_/Q _4201_/A1 VDD VSS
+ gf180mcu_fd_sc_mcu7t5v0__aoi222_1
XTAP_1205 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_70_602 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7958_ _7958_/D _7959_/RN _7958_/CLK _7958_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XTAP_1238 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1227 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1216 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_70_613 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7889_ _7889_/D _7901_/RN _7889_/CLK _7889_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffsnq_1
XTAP_1249 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_23_540 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_23_551 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_24_11 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6909_ _6953_/A2 _6941_/A2 _6908_/Z _7194_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor3_4
XFILLER_168_534 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_23_562 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_50_392 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_155_239 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_149_792 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_6_205 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_40_32 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_163_283 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_151_445 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_151_423 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_108_199 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_6_2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xhold290 hold290/I _7852_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
XFILLER_78_724 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_77_212 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_46_632 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_65_73 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_46_676 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_18_389 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1761 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1750 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_61_657 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_14_540 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1783 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1794 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1772 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_159_567 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_146_206 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_139_291 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_127_420 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_154_250 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_182_592 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_170_743 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_114_114 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_5240_ _5385_/B2 _5687_/B _5690_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_2
XFILLER_142_467 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5171_ _5171_/A1 _5171_/A2 _5171_/A3 _5171_/A4 _5191_/B1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand4_1
XFILLER_69_724 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_39_2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4122_ hold118/Z _3869_/I _4883_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_4053_ _7761_/Q _6248_/A1 _6384_/A1 _7825_/Q _7841_/Q _6418_/A1 _4057_/A1 VDD VSS
+ gf180mcu_fd_sc_mcu7t5v0__aoi222_1
XFILLER_83_215 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
Xclkbuf_3_0__f_csclk clkbuf_0_csclk/Z _7558_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
Xinput3 debug_out input3/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_49_492 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_92_760 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_64_451 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_37_676 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7812_ _7812_/D _7901_/RN _7812_/CLK _7812_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_64_473 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4955_ _4943_/Z _4955_/A2 _4957_/A4 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_7743_ _7743_/D _7901_/RN _7743_/CLK _7743_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_51_123 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3906_ _3906_/A1 _3906_/A2 _3906_/A3 _3906_/A4 _3917_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand4_1
X_7674_ _7674_/D _7961_/RN _7689_/CLK _7674_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
X_4886_ hold572/Z _4887_/A2 _4887_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_32_392 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_137_206 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3837_ _4153_/A1 hold146/Z _6022_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_4
X_6625_ _7432_/D _6625_/A2 _6625_/B _7920_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_165_559 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_3768_ _7969_/Q _7970_/Q _3772_/S _7970_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_118_442 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6556_ _7435_/Q _7433_/Q _6556_/B _6557_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_173_570 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5507_ _5648_/A1 _5793_/A2 _5624_/B _5648_/B2 _5649_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_106_615 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_161_721 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_145_283 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3699_ _7711_/Q _3699_/ZN VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_105_114 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6487_ hold765/Z _6502_/A2 _6488_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_133_478 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_126_24 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5438_ _5721_/B _5424_/Z _5438_/A3 _5439_/A4 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor3_1
Xoutput340 _7503_/Q wb_dat_o[7] VDD VSS gf180mcu_fd_sc_mcu7t5v0__buf_8
X_5369_ _3728_/I _4996_/Z _5369_/B _5370_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_114_670 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_99_370 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_86_28 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_59_212 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7108_ _7433_/Q _7935_/Q _7106_/Z _7108_/B2 _7109_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_7039_ _7035_/Z _7039_/A2 _7039_/A3 _7039_/A4 _7054_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand4_1
XFILLER_75_705 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_75_716 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_28_676 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1002 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1013 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1035 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1046 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1024 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_43_668 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_70_487 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1079 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1068 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1057 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_156 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_168_353 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_143_2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_136_250 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_136_272 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_151_242 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_3_753 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_808 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_151_286 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_2_274 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_819 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_120_673 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_76_61 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_65_215 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_19_632 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_34_602 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_46_495 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_2270 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_73_292 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_18_197 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2292 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2281 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_92_93 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4740_ hold562/Z _4740_/I1 _4741_/S _4740_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XTAP_1591 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1580 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_14_392 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_42_690 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4671_ hold55/I hold41/Z hold42/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_174_323 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_147_559 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6410_ hold392/Z _6417_/A2 _6411_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_7390_ _7390_/D _7961_/RN _7874_/CLK _7390_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
X_6341_ hold73/Z _6349_/A2 _6341_/B _7801_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_155_570 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_127_283 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_115_412 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_170_540 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6272_ hold373/Z _6281_/A2 _6273_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_5223_ _5302_/A1 _5195_/B _5224_/A3 _5224_/A4 _5433_/C VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor4_4
XFILLER_88_318 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5154_ _5496_/A1 _5543_/B _5153_/C _5552_/A3 _5155_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor4_2
X_4105_ _4105_/A1 _4105_/A2 _4106_/A4 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_84_502 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_5085_ _5496_/A1 _5319_/C _5660_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_4036_ _4025_/Z _4036_/A2 _4036_/A3 _4036_/A4 _4036_/ZN VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor4_1
XFILLER_112_37 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_107 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
X_5987_ hold90/Z _5987_/A2 _5987_/B hold222/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
XPHY_129 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_118 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_12_318 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_40_605 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7726_ _7726_/D _7901_/RN _7755_/CLK _7726_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffsnq_1
X_4938_ _4941_/C _4941_/B _4942_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_178_673 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7657_ _7657_/D _7961_/RN _7735_/CLK _7657_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
X_4869_ hold687/Z _4872_/A2 _4870_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_6608_ _6586_/B _6608_/A2 _6611_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_153_507 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_137_12 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_118_250 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7588_ _7588_/D input75/Z _7589_/CLK _7998_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_134_721 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6539_ _4448_/Z _6553_/A2 _6539_/B _7894_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_137_67 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_134_743 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_106_467 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_133_275 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_133_286 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_121_404 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
Xoutput170 _4433_/Z irq[2] VDD VSS gf180mcu_fd_sc_mcu7t5v0__buf_8
Xoutput181 _3693_/ZN mgmt_gpio_oeb[19] VDD VSS gf180mcu_fd_sc_mcu7t5v0__buf_8
Xoutput192 _3683_/ZN mgmt_gpio_oeb[29] VDD VSS gf180mcu_fd_sc_mcu7t5v0__buf_8
XFILLER_102_673 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_47_204 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_75_546 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_47_215 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_56_760 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_46_53 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_46_86 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XPHY_9 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_43_421 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_55_281 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_71_774 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_71_785 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_102_92 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_62_41 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_31_638 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_8_812 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_7_311 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_137_570 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_109_283 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_171_348 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_98_605 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_605 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_616 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_140_768 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_627 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_638 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_649 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_78_362 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_66_524 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5910_ hold167/Z hold276/I _5911_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_6890_ _7475_/Q _6890_/A2 _6890_/B1 _7396_/Q _6896_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_46_270 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_61_240 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5841_ _5841_/A1 _7285_/A2 _5845_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_22_605 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_5772_ _5772_/A1 _5173_/B _5772_/A3 _5773_/C VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand3_1
X_7511_ _7511_/D _7959_/RN _7958_/CLK _7511_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffsnq_1
X_4723_ _4454_/Z _4731_/A2 _4723_/B _7445_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_7442_ hold87/Z _7961_/RN _7603_/CLK _7442_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_30_671 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_175_665 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4654_ _7424_/Q _4685_/A1 _4657_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_1
Xinput61 mgmt_gpio_in[32] input61/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
Xinput50 mgmt_gpio_in[22] input50/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
Xinput72 mgmt_gpio_in[9] input72/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_7373_ _7373_/D _7901_/RN _7876_/CLK _7373_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
X_4585_ hold648/Z _4588_/A2 _4586_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_162_348 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_143_540 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6324_ hold73/Z _6332_/A2 _6324_/B _7793_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
Xinput83 spimemio_flash_clk input83/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
Xinput94 uart_enabled _4400_/S VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_131_702 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6255_ hold531/Z _6264_/A2 _6256_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_89_638 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_88_104 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_170_392 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5206_ _5369_/B _5206_/A2 _5205_/Z _5207_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor3_1
XFILLER_115_286 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6186_ hold283/Z _6191_/A2 _6187_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_88_159 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_5137_ _5309_/A1 _3723_/I _5344_/A1 _5498_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand3_4
XFILLER_123_25 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_96_181 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_96_170 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_84_321 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_29_215 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5068_ _5302_/A1 _5211_/A3 _4920_/Z _5069_/A4 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand3_2
XFILLER_29_237 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_83_29 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4019_ _7656_/Q _6022_/A1 _5971_/A1 _7632_/Q _4020_/A4 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_72_527 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_65_590 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_16_34 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_37_270 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_80_582 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_80_593 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_13_638 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7709_ _7709_/D _7901_/RN _7812_/CLK _7709_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffsnq_1
XFILLER_8_108 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_32_33 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_32_55 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_166_676 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_148_33 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_21_693 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_138_389 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_126_529 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_119_570 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_107_721 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_106_2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_180_189 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_180_167 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_79_115 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_164_76 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_122_735 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_121_212 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_76_811 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_597 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_48_513 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_75_354 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_48_568 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_63_549 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_73_73 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_16_454 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_71_593 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_43_273 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_172_602 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_7_141 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_156_164 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xhold108 hold108/I hold108/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
X_4370_ _4924_/A3 _4924_/A4 _4370_/A3 _4370_/A4 _4372_/A4 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor4_1
XFILLER_172_657 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
Xhold119 hold119/I hold119/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
XFILLER_152_392 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_98_446 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_424 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_402 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_413 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_6040_ hold673/Z _6055_/A2 _6041_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_112_256 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_457 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_446 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_435 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_66_321 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_479 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_468 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_21_2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_93_140 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_66_343 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7991_ _7991_/I _7991_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_94_696 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6942_ _7189_/A2 _7191_/A2 _7197_/A2 _7193_/B1 _6946_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor4_1
XFILLER_81_357 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_62_560 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6873_ _6873_/A1 _6867_/Z _6873_/A3 _6875_/B1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand3_1
X_5824_ hold495/Z _5827_/A2 _5825_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_35_785 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_50_744 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_22_457 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5755_ _5755_/A1 _5755_/A2 _5777_/B _5756_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi21_1
Xclkbuf_leaf_90_csclk _7558_/CLK _7875_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_148_676 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4706_ _4718_/A1 hold173/Z _4706_/B hold174/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_5686_ _5363_/B _5686_/A2 _5627_/Z _5686_/A4 _5686_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__and4_1
XFILLER_163_635 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4637_ _7994_/I _4652_/A1 _4640_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_7425_ hold38/Z _7901_/RN _7816_/CLK _7425_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_147_175 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
Xhold620 _7410_/Q hold620/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
Xhold642 _7806_/Q hold642/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
XFILLER_150_318 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xhold653 _7585_/Q hold653/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
XFILLER_78_29 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_7356_ _7356_/D _7961_/RN _7370_/CLK _7356_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffsnq_2
XFILLER_1_306 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xhold631 _7637_/Q hold631/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
X_4568_ _4454_/Z _4568_/A2 _4568_/B _7390_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
Xhold675 _7724_/Q hold675/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
XFILLER_103_201 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_103_212 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_103_223 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6307_ hold73/Z _6315_/A2 _6307_/B _7785_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_4499_ hold539/Z _4504_/A2 hold540/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
Xhold686 _7538_/Q hold686/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
X_7287_ _4448_/Z _7289_/A2 _7287_/B _7960_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
Xhold697 _7393_/Q hold697/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
Xhold664 _7407_/Q hold664/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
X_6238_ hold47/Z _6242_/A2 _6238_/B _7753_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_89_457 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6169_ hold422/Z _6174_/A2 _6170_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_980 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_134_79 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_85_641 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_991 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_57_387 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
Xclkbuf_leaf_43_csclk clkbuf_3_7__f_csclk/Z _7461_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_150_34 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_57_398 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_13_413 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_53_582 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_25_295 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_159_65 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xclkbuf_leaf_58_csclk _7961_/CLK _7815_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_9_428 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_40_254 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_43_98 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_138_131 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_127_805 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_166_473 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_138_164 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_5_623 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_181_432 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_175_53 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_154_646 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_5_645 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_5_634 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_4_133 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_134_392 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_4_188 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_4_37 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_108_91 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_48_321 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_124_90 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_75_140 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_63_357 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_90_176 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_17_785 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_32_711 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_176_204 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3870_ _4075_/B _3869_/I _4505_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_4
XFILLER_176_259 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_290 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
X_5540_ _5735_/A2 _5179_/B _5540_/B1 _5540_/B2 _5540_/C _5642_/A4 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi221_2
XFILLER_172_410 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5471_ _5674_/A1 _5471_/A2 _5749_/A3 _5471_/A4 _5472_/C VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand4_1
XFILLER_8_472 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_69_2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4422_ _4422_/I _4422_/ZN VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_7210_ _7210_/A1 _7210_/A2 _7210_/B _7433_/Q _7211_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XFILLER_160_605 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_132_318 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_160_649 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_132_329 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7141_ _7877_/Q _7195_/C1 _7193_/C1 _7731_/Q _7667_/Q _7194_/B1 _7144_/A2 VDD VSS
+ gf180mcu_fd_sc_mcu7t5v0__aoi222_1
X_4353_ _6905_/A1 _7916_/Q _6937_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_4
XFILLER_101_716 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_99_766 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_7072_ _7826_/Q _7202_/A2 _7204_/B1 _7770_/Q _7077_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_4284_ _4284_/A1 _4427_/B _7219_/A1 _4284_/B _7548_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai31_1
XFILLER_99_799 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6023_ hold768/Z _6038_/A2 _6024_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_104_27 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_67_641 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7974_ _7974_/D _7327_/Z _7977_/CLK _7974_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_67_696 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1409 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_81_154 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6925_ _7912_/Q _7911_/Q _6936_/A2 _6951_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand3_4
XFILLER_120_37 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_168_727 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_6856_ _7529_/Q _6881_/A2 _6881_/B1 _7523_/Q _6859_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_167_215 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6787_ _6787_/A1 _6787_/A2 _6787_/A3 _6792_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand3_1
X_3999_ _3999_/A1 _3999_/A2 _3999_/A3 _3998_/Z _7227_/I0 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand4_4
XFILLER_10_405 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5807_ _5807_/A1 _7285_/A2 _5811_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_148_451 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5738_ _5698_/B _5738_/A2 _5738_/B _5738_/C _5756_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_136_646 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_5669_ _5669_/A1 _5179_/B _5669_/B _5799_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_108_337 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_89_28 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_123_318 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7408_ _7408_/D _7961_/RN _7756_/CLK _7408_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
X_7339_ _7339_/D _7294_/Z _4415_/A2 _7339_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_151_638 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xhold472 _7851_/Q hold472/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
Xhold461 _7772_/Q hold461/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
XFILLER_116_392 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xhold450 _7837_/Q hold450/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
XFILLER_89_210 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_8_6 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_150_148 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_145_67 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xhold483 _7562_/Q hold483/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
Xhold494 _7447_/Q hold494/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
XFILLER_85_460 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_38_65 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_45_302 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_173_2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_161_99 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_18_538 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1910 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_45_357 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1943 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1932 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1921 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1976 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1965 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1954 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_14_744 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1998 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1987 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_139_473 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_70_74 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_182_752 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_126_134 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_181_240 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_142_605 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_114_318 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_79_61 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_79_50 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_96_747 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_96_769 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_96_758 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_68_449 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_49_630 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_49_641 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_49_663 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_91_463 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_52_806 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4971_ _5006_/B _5254_/A2 _5206_/A2 _5104_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor3_4
XFILLER_91_496 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_91_474 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_7690_ _7690_/D _7961_/RN _7691_/CLK _7690_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
X_6710_ _7133_/S _6710_/A2 _6710_/B _7922_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_3922_ _4402_/A1 _4427_/B _3922_/B _7555_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_32_530 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_149_226 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_149_215 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3853_ _4212_/A2 hold133/Z _6452_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_4
X_6641_ _7910_/Q _6663_/A4 _6658_/A3 _6885_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor3_4
XFILLER_165_708 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_20_747 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_158_771 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3784_ _3810_/S hold122/Z _3784_/B hold123/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi21_4
XFILLER_118_624 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_118_602 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6572_ _6572_/A1 _4352_/B _6618_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_2
X_5523_ _5519_/B _5559_/A1 _5523_/A3 _5524_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__or3_1
X_5454_ _5783_/A2 _5668_/A2 _5454_/B _5460_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_117_156 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5385_ _5603_/A1 _4993_/B _4993_/C _5409_/B2 _5385_/B2 _5583_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai32_1
X_4405_ _7424_/Q input3/Z input1/Z _4405_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_7124_ _7884_/Q _7203_/B1 _7204_/A2 _7844_/Q _7129_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_4336_ _7978_/Q hold11/I _4338_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_87_703 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_115_15 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7055_ _7607_/Q _7210_/A2 _7055_/B _7433_/Q _7058_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi211_1
X_4267_ _4267_/A1 _4267_/A2 _4267_/A3 _4267_/A4 _4281_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand4_1
X_6006_ hold772/Z _6021_/A2 _6007_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_4198_ _4198_/A1 _4198_/A2 _4198_/A3 _4198_/A4 _4202_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand4_1
XFILLER_95_780 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_82_463 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_15_508 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_27_357 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7957_ _7957_/D _7959_/RN _4411_/I1 hold88/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_131_69 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1239 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1228 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1217 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1206 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_7888_ _7888_/D _7901_/RN _7893_/CLK _7888_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
X_6908_ _6908_/A1 _7913_/Q _6908_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__or2_4
X_6839_ _6839_/A1 _6839_/A2 _6839_/A3 _6848_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_24_45 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_24_34 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_7_707 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_108_101 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_7_718 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_164_752 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_156_33 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_124_605 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_156_77 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
Xhold280 _7714_/Q hold280/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
XFILLER_172_21 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
Xhold291 _7712_/Q hold291/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
XFILLER_78_747 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_77_235 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_49_97 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_58_460 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_65_85 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_61_603 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_45_176 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1751 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1740 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1784 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1773 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1762 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_60_179 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_147_708 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1795 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_81_73 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_155_785 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_142_402 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_127_476 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_115_638 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_6_784 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_142_457 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_5_283 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5170_ _5666_/A1 _5658_/B _5179_/B _5672_/A2 _5171_/A4 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_110_321 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_96_555 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_96_544 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_68_235 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_4121_ hold133/Z hold107/Z _4589_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_110_376 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_96_566 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4052_ _4052_/A1 _4052_/A2 _4052_/A3 _4058_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand3_1
Xinput4 mask_rev_in[0] input4/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_37_633 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_7811_ _7811_/D _7901_/RN _7812_/CLK _7811_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_64_463 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_36_165 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_51_102 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4954_ _5069_/A2 _4930_/Z _4953_/Z _5661_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand3_4
X_7742_ _7742_/D _7901_/RN _7849_/CLK _7742_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffsnq_1
XFILLER_52_647 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3905_ input60/Z _5886_/A1 _6537_/A1 _7901_/Q _3906_/A4 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_177_354 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7673_ _7673_/D _7901_/RN _7673_/CLK _7673_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_60_680 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4885_ _4448_/Z _4887_/A2 _4885_/B _7533_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_3836_ _4153_/A1 _3835_/Z _5937_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_4
X_6624_ _7920_/Q _6625_/A2 _6625_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_3767_ _7970_/Q _7971_/Q _3772_/S _7971_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_6555_ _7435_/Q _7433_/Q _6562_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_161_700 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5506_ _5735_/A2 _5179_/B _5540_/C _5506_/C _5508_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XFILLER_106_605 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_145_295 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3698_ _7719_/Q _3698_/ZN VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_6486_ _6486_/A1 _7285_/A2 _6502_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_4
X_5437_ _5714_/B1 _5722_/A1 _5437_/B _5438_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
Xoutput330 _7945_/Q wb_dat_o[27] VDD VSS gf180mcu_fd_sc_mcu7t5v0__buf_8
Xoutput341 _7486_/Q wb_dat_o[8] VDD VSS gf180mcu_fd_sc_mcu7t5v0__buf_8
X_5368_ _5689_/A1 _5618_/B1 _5565_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_161_799 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_126_69 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_114_660 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_102_811 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_86_18 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5299_ _5173_/C _5299_/A2 _5299_/A3 _5299_/A4 _5300_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand4_1
X_4319_ _4309_/S _4319_/A2 _4319_/B _7338_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_113_181 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_7107_ _7107_/A1 _7210_/A2 _7433_/Q _7108_/B2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_59_224 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_101_354 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7038_ _7817_/Q _7207_/A2 _7205_/B1 _7743_/Q _7039_/A4 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_47_419 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_142_46 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_74_238 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_83_783 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_35_22 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_43_625 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1003 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_169_800 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1036 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1047 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1025 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_35_55 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_55_496 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1014 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_168_321 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_70_477 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1069 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1058 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_179 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_70_499 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_156_527 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_136_2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_11_566 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_156_538 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_51_65 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_137_763 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_109_443 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_137_785 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_152_755 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_152_744 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_111_107 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_809 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_104_170 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_78_555 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_78_544 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_65_227 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_19_611 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_81_709 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_74_761 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_18_176 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_46_463 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_2271 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2260 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_73_282 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2293 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2282 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_159_354 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1592 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1581 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1570 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_61_499 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_42_680 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4670_ _7985_/I _4685_/A1 _4673_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_174_335 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_6340_ hold496/Z _6349_/A2 _6341_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_51_2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6271_ _4460_/Z _6281_/A2 _6271_/B _7768_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_5222_ _5376_/B _5392_/B2 _5294_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_115_479 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5153_ _5552_/A3 _5539_/A3 _5543_/B _5153_/C _5180_/C1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XFILLER_111_641 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4104_ _4104_/A1 _4104_/A2 _4104_/A3 _4104_/A4 _4105_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand4_1
X_5084_ _5643_/A2 _5087_/B _5600_/B2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_110_173 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_110_195 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_4035_ _4035_/A1 _4035_/A2 _4035_/A3 _4035_/A4 _4036_/A4 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand4_1
XFILLER_65_783 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_64_260 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_37_463 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_37_496 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_52_444 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5986_ hold221/Z _5987_/A2 _5987_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XPHY_119 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_52_455 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_108 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
X_4937_ _5200_/B _3727_/I _4946_/A1 _5230_/A1 _4941_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor4_4
X_7725_ _7725_/D _7901_/RN _7753_/CLK _7725_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffsnq_1
XFILLER_24_179 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_52_499 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_177_140 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7656_ _7656_/D _7961_/RN _7702_/CLK _7656_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
X_4868_ _4868_/A1 _7285_/A2 _4872_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_3819_ hold630/I _3817_/I _3819_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__or2_4
X_6607_ _7434_/Q _6610_/A3 _6608_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_180_305 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_165_357 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7587_ _7587_/D _7961_/RN _7587_/CLK _7587_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
X_4799_ _7486_/Q _4809_/S _4800_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_119_785 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_115_7 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6538_ hold738/Z _6553_/A2 _6539_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_134_755 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6469_ _6469_/A1 _7285_/A2 _6485_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_4
XFILLER_0_702 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_153_12 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_99_190 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
Xoutput171 _4409_/ZN mgmt_gpio_oeb[0] VDD VSS gf180mcu_fd_sc_mcu7t5v0__buf_8
Xoutput182 _4407_/ZN mgmt_gpio_oeb[1] VDD VSS gf180mcu_fd_sc_mcu7t5v0__buf_8
Xoutput193 _3710_/ZN mgmt_gpio_oeb[2] VDD VSS gf180mcu_fd_sc_mcu7t5v0__buf_8
XFILLER_75_503 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_768 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_101_173 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_75_514 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_101_184 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_63_709 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_46_32 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_90_517 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_28_463 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_55_271 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_70_241 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_15_168 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_169_641 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_30_105 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_43_499 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_11_374 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_144_519 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_97_105 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_3_540 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_606 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_140_747 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_112_427 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_97_138 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_617 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_628 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_639 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_94_812 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_120_460 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_66_514 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_46_260 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_47_783 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_19_496 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5840_ hold47/Z _5840_/A2 _5840_/B _7568_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_34_444 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_34_477 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_2090 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_5771_ _5771_/A1 _5805_/A1 _5805_/B _5787_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_99_2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4722_ hold635/Z _4731_/A2 _4723_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_7510_ _7510_/D _7961_/RN _7510_/CLK _7510_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
X_7441_ hold59/Z _7901_/RN _7583_/CLK _7441_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_174_121 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_159_184 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_147_357 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4653_ _4653_/A1 _5903_/A2 _4686_/B1 hold55/Z hold12/Z _4685_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi221_4
Xinput40 mgmt_gpio_in[13] input40/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_174_176 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xinput62 mgmt_gpio_in[33] input62/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
Xinput51 mgmt_gpio_in[23] input51/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
Xinput73 pad_flash_io0_di input73/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_7372_ _7372_/D _7901_/RN _7573_/CLK _7372_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
X_4584_ _4584_/A1 _7285_/A2 _4588_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
Xinput95 wb_adr_i[0] _3723_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__buf_16
X_6323_ hold502/Z _6332_/A2 _6324_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_128_593 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_116_744 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_115_221 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_115_210 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
Xinput84 spimemio_flash_csb input84/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_6254_ _4460_/Z _6264_/A2 _6254_/B hold262/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_5205_ _5338_/A1 _4996_/Z _5205_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_130_213 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_103_449 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6185_ hold41/Z _6191_/A2 _6185_/B _7728_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_85_812 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5136_ _5136_/A1 _5344_/A2 _5680_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_2
XFILLER_123_15 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5067_ _3722_/I _5087_/C _5344_/A1 _5527_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand3_4
XFILLER_84_333 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_45_709 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4018_ input24/Z _4239_/A2 _6282_/A1 _7778_/Q _4020_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_53_742 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_80_550 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_16_68 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_25_444 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_80_572 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_12_105 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5969_ hold308/Z _5970_/A2 _5970_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_25_499 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7708_ _7708_/D _7901_/RN _7812_/CLK _7708_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffsnq_1
XFILLER_178_471 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_32_45 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_148_56 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7639_ _7639_/D _7961_/RN _7645_/CLK _7639_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_166_699 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_165_176 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_153_316 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_180_179 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_106_254 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_122_747 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_94_108 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_554 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_102_460 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_87_171 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_180_65 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_29_783 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_63_539 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_56_591 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_73_96 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_31_425 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_129_357 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_11_171 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_11_160 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_8_654 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_156_187 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_156_176 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_129_379 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_8_676 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_171_124 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xhold109 hold109/I _7446_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
XFILLER_171_179 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_125_552 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_113_736 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_98_436 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_98_425 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_3_370 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_403 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_414 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_98_458 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_458 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_447 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_436 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_425 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_121_780 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_67_812 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_469 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_82_804 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_14_2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_27_709 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7990_ _7990_/I _7990_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_94_686 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_6941_ _6941_/A1 _6941_/A2 _7196_/B1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_4
XFILLER_34_230 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_35_775 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6872_ _7525_/Q _6889_/A2 _6853_/Z _6830_/B _6872_/C _6873_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi221_1
XFILLER_62_572 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5823_ _4460_/Z _5827_/A2 _5823_/B _7560_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_5754_ _5754_/A1 _5754_/A2 _5754_/A3 _5800_/A1 _5755_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor4_1
X_4705_ hold172/Z _3819_/Z _4705_/B hold173/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_5685_ _5759_/A1 _5724_/A2 _5685_/B _5686_/A4 VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_175_496 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4636_ _4652_/A1 hold83/Z _4636_/B hold84/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_162_102 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_7424_ hold78/Z _7901_/RN _7583_/CLK _7424_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_151_809 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_118_37 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_116_530 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7355_ _7355_/D _7961_/RN _7875_/CLK _7355_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffsnq_1
Xhold621 _7505_/Q hold621/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
Xhold610 _7406_/Q hold610/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
XFILLER_162_179 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_162_157 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xhold643 _7628_/Q hold643/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
X_6306_ hold362/Z _6315_/A2 _6307_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_4567_ hold571/Z _4568_/A2 _4568_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
Xhold654 _7756_/Q hold654/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
Xhold632 _7386_/Q hold632/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
Xhold676 _7375_/Q hold676/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
XFILLER_143_382 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_116_596 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_104_747 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_89_425 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xhold665 _7998_/I hold665/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
X_4498_ hold41/Z _4504_/A2 _4498_/B hold478/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
Xhold687 _7527_/Q hold687/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
X_7286_ hold757/Z _7289_/A2 _7287_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_6237_ hold285/Z _6242_/A2 _6238_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_131_566 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
Xhold698 _7356_/Q hold698/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
X_6168_ hold41/Z _6174_/A2 _6168_/B _7720_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_76_108 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_58_812 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_970 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_57_300 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5119_ _5476_/B _5689_/A2 _7520_/Q _5519_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
XTAP_981 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_992 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_6099_ hold223/Z _6106_/A2 _6100_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_13_425 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_40_211 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_41_712 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_158_408 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_13_447 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_41_745 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_43_33 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_179_780 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_139_611 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_166_463 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_138_176 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_153_124 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_181_499 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_107_596 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_107_585 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_108_81 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_95_406 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_68_63 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_110_717 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_103_780 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_95_428 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_95_417 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_68_96 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_49_812 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_88_480 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_384 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_91_601 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_75_163 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_48_388 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_91_667 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_44_561 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_44_572 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_177_728 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_32_767 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_169_290 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_291 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_280 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_117_316 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5470_ _4969_/C _4996_/Z _5471_/A4 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_157_496 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_8_484 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4421_ _4424_/A1 input86/Z _4422_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_2
XFILLER_144_179 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_99_712 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7140_ _7140_/A1 _7140_/A2 _7140_/A3 _7140_/A4 _7140_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__and4_1
X_4352_ _7001_/C _4361_/A2 _4352_/B _7433_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_152_190 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_99_778 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7071_ _7762_/Q _7202_/C2 _7202_/B1 _7786_/Q _7077_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_4283_ _4283_/A1 _4283_/A2 _4283_/A3 _4283_/A4 _7219_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor4_4
X_6022_ _6022_/A1 hold32/Z _6038_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_4
XFILLER_100_205 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_98_266 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_58_108 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_67_631 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_39_311 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_82_634 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_7973_ _7973_/D _7326_/Z _7977_/CLK _7973_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_66_174 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_81_144 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6924_ _7912_/Q _7911_/Q _6955_/A4 _6908_/Z _7190_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor4_4
XFILLER_23_712 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_168_717 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6855_ _7531_/Q _6892_/B1 _6880_/B1 _7409_/Q _6867_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_50_531 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5806_ _5806_/A1 _5806_/A2 _5806_/A3 _5806_/A4 _7545_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand4_1
X_6786_ _7697_/Q _6881_/B1 _6880_/B1 _7811_/Q _6787_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_3998_ _3998_/A1 _3998_/A2 _3998_/A3 _3998_/A4 _3998_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__and4_1
XFILLER_23_789 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5737_ _5795_/A2 _5737_/A2 _5785_/A1 _5737_/B _5738_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai31_1
XFILLER_148_463 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5668_ _5783_/A2 _5668_/A2 _5668_/B _5668_/C _5776_/A4 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi211_2
XFILLER_129_69 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7407_ _7407_/D _7961_/RN _7756_/CLK _7407_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
X_5599_ _5599_/A1 _5661_/B _5656_/A2 _5665_/A1 _5599_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__and4_1
X_4619_ _5886_/A1 _5903_/A2 _4686_/B1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_4
XFILLER_2_605 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_163_499 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7338_ _7338_/D _7293_/Z _4031_/C2 _7338_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
Xhold440 _7804_/Q hold440/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
Xhold462 _7885_/Q hold462/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
Xhold451 _7704_/Q hold451/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
X_7269_ _7519_/Q _7269_/A2 _7271_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
Xhold473 _7380_/Q hold473/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
Xhold484 _7771_/Q hold484/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
XFILLER_104_555 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_104_566 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_104_544 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
Xhold495 _7561_/Q hold495/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
XFILLER_77_428 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_58_620 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_38_33 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_38_77 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_57_141 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_57_152 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_85_483 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_72_122 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_72_100 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_38_99 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_166_2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1900 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1933 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1922 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1911 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1977 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1966 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1955 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1944 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_26_594 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1999 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1988 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_9_215 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_9_237 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_167_783 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_167_761 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_127_614 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_181_230 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_139_496 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_154_477 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_126_179 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_79_40 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_5_487 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_79_73 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_96_737 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_181 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_1_682 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_36_336 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_63_144 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4970_ _5006_/B _5206_/A2 _5608_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_4
XFILLER_63_166 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_17_550 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_177_503 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3921_ _7554_/Q _4284_/A1 _3921_/B _4427_/B _3922_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi211_1
X_3852_ _3796_/Z _4075_/B _4239_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_4
XFILLER_32_575 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6640_ _7910_/Q _6658_/A2 _6662_/A3 _6889_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor3_4
XFILLER_81_2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6571_ _6557_/I _6571_/A2 _6570_/Z _6564_/B _6571_/B2 _7905_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai32_1
X_5522_ _5522_/A1 _5520_/C _5522_/B1 _5522_/B2 _7540_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_3783_ hold18/Z _3781_/Z _3810_/S hold19/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_4
XFILLER_117_124 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_145_477 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5453_ _5714_/A1 _5527_/A1 _5668_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_2
X_5384_ _5392_/A1 _5392_/A2 _5376_/B _5405_/B _5392_/B2 _5702_/C VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai32_1
Xclkbuf_leaf_42_csclk clkbuf_3_7__f_csclk/Z _7463_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_145_499 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_132_116 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_132_105 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_117_179 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4404_ _7979_/Q _4425_/A2 _4404_/B _4404_/ZN VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi21_2
X_7123_ _7836_/Q _7203_/A2 _7204_/B1 _7772_/Q _7129_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_99_531 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4335_ _7630_/Q _4335_/A2 _5903_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_4
XFILLER_5_70 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_99_597 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_59_417 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_59_428 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_115_49 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_86_247 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7054_ _7054_/A1 _7054_/A2 _7054_/A3 _7054_/A4 _7055_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__or4_1
X_4266_ _7830_/Q _6401_/A1 _4614_/A1 _7409_/Q _4267_/A4 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_1
Xclkbuf_leaf_57_csclk _7961_/CLK _7791_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
X_6005_ _6005_/A1 _7285_/A2 _6021_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_4
XFILLER_39_152 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_39_141 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_39_130 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4197_ _7895_/Q _6537_/A1 _4594_/A1 _7402_/Q _6243_/A1 _7757_/Q _4198_/A4 VDD VSS
+ gf180mcu_fd_sc_mcu7t5v0__aoi222_1
XFILLER_54_100 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_82_442 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_82_431 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7956_ _7956_/D _7959_/RN _4411_/I1 hold66/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XTAP_1229 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1218 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1207 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_7887_ _7887_/D _7901_/RN _7887_/CLK _7887_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
X_6907_ _6953_/A1 _6599_/Z _6941_/A2 _7195_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor3_4
X_6838_ _7382_/Q _6882_/A2 _6882_/B1 _7659_/Q _6839_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_168_558 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_149_783 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6769_ _7680_/Q _6887_/B1 _6891_/B1 _7672_/Q _6771_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_10_258 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_10_247 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_164_742 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_148_282 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_10_269 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_40_34 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_164_797 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_156_56 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_151_425 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_108_179 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_156_89 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xhold270 hold270/I _6221_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
XFILLER_123_138 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xhold292 _7663_/Q hold292/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
Xhold281 _7633_/Q hold281/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
XFILLER_132_683 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_132_672 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_120_812 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_49_32 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_49_65 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_46_601 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_105_93 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_58_483 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_18_325 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_65_64 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_45_144 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1752 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1741 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1730 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_121_70 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_14_531 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1785 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1774 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1763 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_159_558 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1796 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_14_597 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_41_361 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_182_594 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_127_499 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_130_609 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_123_650 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_111_812 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_69_726 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_96_534 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_68_247 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4120_ hold118/Z _3881_/Z _4863_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_4051_ _7857_/Q _6452_/A1 _6401_/A1 _7833_/Q _7809_/Q _6350_/A1 _4052_/A3 VDD VSS
+ gf180mcu_fd_sc_mcu7t5v0__aoi222_1
Xinput5 mask_rev_in[10] input5/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_7810_ _7810_/D _7901_/RN _7810_/CLK _7810_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_92_751 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_25_807 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4953_ _4906_/Z _5138_/A2 _4953_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__and2_4
XFILLER_91_283 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7741_ _7741_/D _7961_/RN _7791_/CLK _7741_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffsnq_1
XFILLER_51_125 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_178_812 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7672_ _7672_/D _7901_/RN _7818_/CLK _7672_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
X_3904_ input51/Z _4275_/A2 _6469_/A1 _7869_/Q _3906_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_4884_ hold751/Z _4887_/A2 _4885_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_6623_ _7432_/Q _7435_/Q _6623_/B _6625_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_118_400 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3835_ hold19/Z _3787_/Z hold127/Z _3794_/Z _3835_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__or4_4
XFILLER_20_534 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3766_ _7971_/Q _7972_/Q _3772_/S _7972_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_6554_ _7433_/Q _4331_/Z _6556_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_173_561 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5505_ _5155_/B _5505_/A2 _5499_/Z _5505_/A4 _5505_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__or4_1
X_6485_ hold90/Z _6485_/A2 _6485_/B _7869_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_161_712 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_160_200 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_160_211 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3697_ _7727_/Q _3697_/ZN VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_133_425 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5436_ _5731_/B _5287_/B _5439_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_106_617 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_10_37 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_126_37 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_105_138 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xoutput331 _7946_/Q wb_dat_o[28] VDD VSS gf180mcu_fd_sc_mcu7t5v0__buf_8
Xoutput342 _7487_/Q wb_dat_o[9] VDD VSS gf180mcu_fd_sc_mcu7t5v0__buf_8
Xoutput320 _7480_/Q wb_dat_o[18] VDD VSS gf180mcu_fd_sc_mcu7t5v0__buf_8
X_5367_ _5774_/A1 _5669_/A1 _5782_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_120_108 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_4318_ _7337_/Q _7414_/Q _4318_/B _4319_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_113_160 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_7106_ _7210_/A2 _7106_/A2 _7106_/A3 _7106_/A4 _7106_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__or4_1
X_5298_ _5580_/A1 _5298_/A2 _5298_/A3 _5298_/A4 _5299_/A4 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor4_1
XFILLER_87_567 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7037_ _7679_/Q _7191_/A2 _7194_/B1 _7663_/Q _7039_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_4249_ input4/Z _4249_/A2 _4764_/A1 _7470_/Q _4253_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_142_25 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_27_144 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_28_656 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_55_420 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_83_795 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_82_250 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_55_475 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_55_486 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_1004 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1037 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1026 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_27_199 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_7939_ _7939_/D _7961_/RN _7940_/CLK _7939_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XTAP_1015 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_169_812 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_70_456 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1059 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1048 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_129_709 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_70_489 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_167_44 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_129_2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_7_538 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_171_509 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_164_594 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_109_499 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_124_458 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_78_534 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_18_100 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_74_751 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_19_689 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_2261 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2250 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_18_188 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_178_108 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2294 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2283 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2272 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_159_311 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1560 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1593 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1582 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1571 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_128_720 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_174_347 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_143_712 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_170_531 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_142_211 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6270_ hold325/Z _6281_/A2 _6271_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_6_582 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5221_ _5585_/A1 _5421_/A1 _5203_/I _5392_/B2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand3_2
XFILLER_142_255 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_102_108 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_44_2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5152_ _5528_/A2 _5020_/Z _5122_/Z _5150_/Z _5546_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand4_2
X_4103_ _7872_/Q _6486_/A1 _6299_/A1 _7784_/Q _6265_/A1 _7768_/Q _4104_/A4 VDD VSS
+ gf180mcu_fd_sc_mcu7t5v0__aoi222_1
XFILLER_57_718 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5083_ _5087_/B _5779_/A1 _5692_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_96_386 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_84_526 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_2_60 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4034_ _7850_/Q _6435_/A1 _5988_/A1 _7640_/Q hold26/I _7575_/Q _4035_/A4 VDD VSS
+ gf180mcu_fd_sc_mcu7t5v0__aoi222_1
XFILLER_64_250 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_24_103 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7724_ _7724_/D _7901_/RN _7813_/CLK _7724_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffsnq_1
X_5985_ hold68/Z _5987_/A2 _5985_/B hold279/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
XPHY_109 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
X_4936_ _5199_/B _5201_/B _4915_/Z _5385_/B2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_165_303 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_138_517 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_7655_ _7655_/D _7961_/RN _7706_/CLK _7655_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
X_4867_ _4454_/Z _4867_/A2 _4867_/B _7526_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_3818_ hold275/Z _3817_/I _5903_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_4
X_7586_ _7586_/D _7961_/RN _7871_/CLK _7586_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
X_6606_ _6953_/A2 _6950_/A2 _6610_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_119_753 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_4798_ _7513_/Q _7959_/RN _4809_/S VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_4
X_6537_ _6537_/A1 _7285_/A2 _6553_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_4
XFILLER_180_328 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_137_36 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_118_252 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_21_69 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3749_ input58/Z _7976_/Q _3749_/S _7976_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_146_594 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_137_58 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_133_233 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_97_29 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_6468_ hold90/Z _6468_/A2 _6468_/B _7861_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_133_277 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5419_ _5087_/B _5292_/B _5419_/B _5419_/C _5727_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi211_2
X_6399_ hold407/Z _6400_/A2 _6400_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_121_406 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xoutput194 _3682_/ZN mgmt_gpio_oeb[30] VDD VSS gf180mcu_fd_sc_mcu7t5v0__buf_8
XFILLER_121_428 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xoutput172 _3702_/ZN mgmt_gpio_oeb[10] VDD VSS gf180mcu_fd_sc_mcu7t5v0__buf_8
Xoutput183 _3692_/ZN mgmt_gpio_oeb[20] VDD VSS gf180mcu_fd_sc_mcu7t5v0__buf_8
XFILLER_0_725 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_153_46 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_101_141 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_153_68 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_47_239 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_56_740 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_83_570 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_46_77 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_15_103 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_55_283 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_62_32 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_43_489 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_178_65 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_7_313 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_7_357 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_137_561 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_125_712 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_124_266 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_607 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_618 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_629 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_87_73 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_87_84 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_39_729 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_93_345 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_16_6 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_46_250 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_53_209 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_179_428 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_61_242 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_61_231 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_34_456 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_34_467 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2091 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2080 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_5770_ _5770_/I _5805_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_61_286 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1390 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_4721_ _4448_/Z _4731_/A2 _4721_/B _7444_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_175_623 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_159_196 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4652_ _4652_/A1 _4652_/A2 _4652_/B hold206/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_7440_ _7440_/D _7961_/RN _7673_/CLK _7989_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_30_673 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xinput30 mask_rev_in[4] input30/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_162_317 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
Xinput63 mgmt_gpio_in[34] input63/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
Xinput41 mgmt_gpio_in[14] input41/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
Xinput52 mgmt_gpio_in[24] input52/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_4583_ _4454_/Z _4583_/A2 _4583_/B _7396_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_7371_ _7371_/D input75/Z _7573_/CLK _7371_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
Xinput96 wb_adr_i[10] input96/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_174_199 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6322_ _4460_/Z _6332_/A2 _6322_/B hold139/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
Xinput85 spimemio_flash_io0_do input85/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
Xinput74 pad_flash_io1_di _3664_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_6253_ hold260/Z _6264_/A2 hold261/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_5204_ _5338_/A1 _5663_/A1 _5381_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_130_203 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_103_428 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6184_ hold329/Z _6191_/A2 _6185_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_130_247 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_97_651 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5135_ _5643_/A2 _5783_/A2 _5765_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_5066_ _5254_/A2 _5448_/A1 _5066_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_84_323 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_29_239 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_57_537 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_84_389 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4017_ _7616_/Q _5937_/A1 _4219_/A2 input16/Z hold114/I _7379_/Q _4020_/A2 VDD VSS
+ gf180mcu_fd_sc_mcu7t5v0__aoi222_1
XFILLER_65_570 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_25_423 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_37_283 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_53_732 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_80_540 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5968_ hold68/Z _5970_/A2 _5968_/B hold348/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_4919_ _5199_/B _5369_/B _4919_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__and2_2
XFILLER_166_601 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7707_ _7707_/D _7961_/RN _7707_/CLK _7707_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_165_111 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_165_100 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5899_ hold335/Z _5902_/A2 _5900_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_21_651 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_165_144 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_165_122 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7638_ _7638_/D _7961_/RN _7642_/CLK _7638_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffsnq_1
XFILLER_32_57 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_148_68 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_107_712 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7569_ _7569_/D _7961_/RN _7875_/CLK _7569_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffsnq_1
XFILLER_134_531 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_134_542 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_180_169 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_164_34 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_107_767 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_164_56 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_79_139 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_130_770 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_102_450 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_88_673 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_48_526 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_180_33 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_28_250 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_16_412 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_44_743 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_43_264 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_43_286 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_85_9 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_12_673 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_12_684 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_172_615 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_140_534 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_404 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_415 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_112_247 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_448 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_437 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_426 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_459 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_94_654 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_94_676 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_94_665 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6940_ _6950_/A1 _6950_/A2 _6941_/A2 _7207_/B1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor3_4
XFILLER_93_175 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_66_389 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_19_283 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_47_570 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_81_359 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6871_ _6871_/A1 _6871_/A2 _6871_/A3 _6872_/C VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand3_1
X_5822_ hold241/Z _5827_/A2 _5823_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_34_264 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_148_601 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5753_ _5099_/B _5753_/A2 _5753_/B _5753_/C _5800_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai211_1
X_4704_ _3819_/Z hold41/Z _4705_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_147_144 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5684_ _5701_/C _5684_/A2 _5684_/A3 _5684_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__and3_1
X_4635_ hold82/Z _3830_/Z _4635_/B hold83/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_7423_ _7423_/D _7901_/RN _7849_/CLK _7997_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
X_7354_ _7354_/D _7961_/RN _7627_/CLK _7354_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffsnq_2
Xhold600 hold600/I _4773_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
X_4566_ _4448_/Z _4568_/A2 _4566_/B _7389_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
Xhold611 _7547_/Q hold611/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
XFILLER_143_350 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6305_ _4460_/Z _6315_/A2 _6305_/B _7784_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
Xhold644 _7759_/Q hold644/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
Xhold633 _7613_/Q hold633/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
Xhold622 hold622/I _4835_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
XFILLER_103_225 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_89_437 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
Xhold688 _7839_/Q hold688/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
Xhold666 _7507_/Q hold666/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
X_4497_ hold476/Z _4504_/A2 hold477/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
Xhold677 _7474_/Q hold677/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
X_7285_ _7285_/A1 _7285_/A2 _7289_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
Xhold655 _7879_/Q hold655/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
X_6236_ hold41/Z _6242_/A2 _6236_/B _7752_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
Xhold699 hold699/I _4492_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
X_6167_ hold327/Z _6174_/A2 _6168_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_134_37 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_112_770 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_960 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_971 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_5118_ _5309_/A1 _3723_/I _4898_/Z _5689_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand3_4
XTAP_982 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_993 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_57_345 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6098_ hold73/Z _6106_/A2 _6098_/B _7687_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_85_687 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_73_805 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_5049_ _5309_/A1 _3723_/I _5006_/B _5448_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor3_4
XFILLER_27_68 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_53_584 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_80_392 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_9_408 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_25_286 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_139_634 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_178_280 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_159_89 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_181_445 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_181_434 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_111_2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_107_531 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_107_520 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_5_625 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_4_113 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_175_77 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_4_135 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_150_810 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_4_179 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_122_534 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_352 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_88_492 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_76_676 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_63_304 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_84_63 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_29_570 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_36_529 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_90_167 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_140_91 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_31_212 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_32_757 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_270 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_292 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_281 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_129_111 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_145_626 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_129_155 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_129_144 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_117_306 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_8_463 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_144_125 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4420_ _4420_/I _4420_/ZN VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_172_467 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4351_ _4331_/Z _6622_/A2 _6569_/A3 _4361_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor3_2
X_7070_ _7882_/Q _7203_/B1 _7204_/A2 _7842_/Q _7834_/Q _7203_/A2 _7077_/A1 VDD VSS
+ gf180mcu_fd_sc_mcu7t5v0__aoi222_1
X_4282_ _4282_/A1 _4282_/A2 _4283_/A4 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_140_375 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_113_567 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6021_ hold90/Z _6021_/A2 _6021_/B hold337/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_67_610 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_82_602 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_39_367 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7972_ _7972_/D _7325_/Z _4415_/A2 _7972_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_94_495 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_82_624 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_67_698 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_54_337 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_54_348 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_54_359 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6923_ _7914_/Q _7913_/Q _6950_/A1 _6955_/A4 _7201_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor4_4
XFILLER_62_392 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6854_ _7401_/Q _6893_/A2 _6890_/B1 _7395_/Q _6867_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_5805_ _5805_/A1 _5804_/Z _5805_/B _5806_/A4 VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_6785_ _7721_/Q _6881_/A2 _6882_/B1 _7657_/Q _6787_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_3997_ _7883_/Q _6503_/A1 _4232_/A2 input8/Z _3997_/C _3998_/A4 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi221_1
XFILLER_22_267 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_23_768 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_23_779 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5736_ _5736_/A1 _5736_/A2 _5706_/Z _5736_/A4 _5785_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand4_2
XFILLER_182_209 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5667_ _5667_/A1 _5602_/Z _5667_/A3 _5748_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_175_283 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_129_59 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_7406_ _7406_/D _7901_/RN _7582_/CLK _7406_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
X_4618_ _4454_/Z _4618_/A2 _4618_/B _7410_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_5598_ _5087_/C _5579_/B _5777_/A2 _5777_/A1 _5665_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_7337_ _7337_/D _7292_/Z _4031_/C2 _7337_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
Xhold463 _7845_/Q hold463/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
XFILLER_89_212 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xhold452 _7696_/Q hold452/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
Xhold441 _7608_/Q hold441/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
X_4549_ _4549_/A1 _7285_/A2 _4553_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
Xhold430 _7353_/Q hold430/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
X_7268_ _7268_/A1 _7277_/B _7268_/B _7955_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi21_1
Xhold485 _7849_/Q hold485/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
Xhold474 _7827_/Q hold474/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
Xhold496 _7801_/Q hold496/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
XFILLER_104_534 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6219_ hold41/Z _6225_/A2 _6219_/B _7744_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_131_364 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_131_353 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_89_267 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_7199_ _7199_/A1 _7199_/A2 _7198_/Z _7209_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_73_602 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_58_676 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_790 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_161_79 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_161_57 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_85_495 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1901 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1934 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1923 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1912 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_72_189 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_60_318 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_54_33 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_159_2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1967 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1956 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1945 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_13_212 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_26_584 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1989 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1978 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_110_50 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_70_32 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_166_250 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_182_787 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_154_467 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_154_456 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_119_81 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_181_286 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_141_117 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_119_92 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_5_499 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_150_673 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_96_727 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_95_215 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_49_621 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_95_73 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_64_602 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_49_665 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_36_315 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_48_175 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_17_540 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3920_ _7976_/Q _7413_/Q _4427_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_4
XFILLER_17_584 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_44_392 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3851_ hold124/Z hold133/Z _6350_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_4
X_3782_ _7506_/Q hold18/Z _3784_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__and2_1
X_6570_ _7905_/Q _6570_/A2 _6570_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_5521_ _5521_/A1 _5521_/A2 _5522_/B2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_74_2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_157_294 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_157_283 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_118_626 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_9_783 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5452_ _4993_/C _5527_/A1 _5543_/C _5452_/C _5454_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XFILLER_173_798 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5383_ _5576_/B2 _5382_/Z _5565_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_4403_ _7334_/Q input38/Z _4403_/B _7979_/Q _4404_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XFILLER_160_459 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7122_ _7828_/Q _7202_/A2 _7202_/B1 _7788_/Q _7764_/Q _7202_/C2 _7129_/A1 VDD VSS
+ gf180mcu_fd_sc_mcu7t5v0__aoi222_1
X_4334_ _7630_/Q _4335_/A2 _4334_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__and2_4
XFILLER_5_82 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_141_684 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_7053_ _7053_/A1 _7053_/A2 _7053_/A3 _7053_/A4 _7054_/A4 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand4_1
XFILLER_101_526 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6004_ hold90/Z _6004_/A2 _6004_/B hold312/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_4265_ _7569_/Q _5841_/A1 _4599_/A1 _7403_/Q _4267_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_4196_ _7557_/Q _5812_/A1 _4754_/A1 _7467_/Q _4198_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_67_495 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_27_348 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_55_646 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7955_ _7955_/D _7959_/RN _4411_/I1 hold45/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XTAP_1219 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1208 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_70_605 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_42_318 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_54_156 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6906_ _6599_/Z _6950_/A2 _6941_/A2 _7189_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor3_4
X_7886_ _7886_/D input75/Z _7886_/CLK _7886_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffsnq_1
X_6837_ _7723_/Q _6881_/A2 _6881_/B1 _7699_/Q _6839_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_148_250 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6768_ _7624_/Q _6659_/Z _6884_/B1 _7688_/Q _6771_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_7_709 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5719_ _5719_/A1 _5677_/Z _5719_/A3 _5719_/A4 _7542_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__or4_1
X_6699_ _7645_/Q _6880_/C2 _6881_/B1 _7693_/Q _7807_/Q _6880_/B1 _6702_/A1 VDD VSS
+ gf180mcu_fd_sc_mcu7t5v0__aoi222_1
XFILLER_163_242 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_124_607 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_108_158 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_163_286 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_108_169 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
Xhold271 hold271/I _7745_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
Xhold260 _7760_/Q hold260/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
XFILLER_104_331 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xhold293 hold293/I _6047_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
Xhold282 hold282/I _7633_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
XFILLER_132_662 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_172_34 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_172_45 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_77_215 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_172_67 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_105_83 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_65_32 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_18_315 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_73_443 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_73_421 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_73_432 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_58_495 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_60_104 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1742 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1731 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1720 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_61_638 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_26_392 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1775 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1764 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1753 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_121_93 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_159_548 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1797 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1786 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_167_570 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_139_283 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_182_562 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_182_551 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_127_467 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_154_275 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_5_241 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_107_191 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_69_705 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_110_334 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4050_ _7873_/Q _6486_/A1 _6039_/A1 _7663_/Q _6022_/A1 _7655_/Q _4052_/A2 VDD VSS
+ gf180mcu_fd_sc_mcu7t5v0__aoi222_1
XFILLER_49_451 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_110_389 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xinput6 mask_rev_in[11] input6/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_92_730 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_36_112 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_24_318 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_52_605 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4952_ _5496_/A1 _5741_/A1 _5602_/A1 _7518_/Q _5474_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai31_1
X_7740_ _7740_/D _7901_/RN _7810_/CLK _7740_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffsnq_1
X_3903_ _7877_/Q _6486_/A1 _6005_/A1 _7651_/Q _6520_/A1 _7893_/Q _3906_/A2 VDD VSS
+ gf180mcu_fd_sc_mcu7t5v0__aoi222_1
X_7671_ _7671_/D _7961_/RN _7735_/CLK _7671_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
X_4883_ _4883_/A1 _7285_/A2 _4887_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_3834_ hold275/Z hold146/Z _5886_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_4
XFILLER_60_682 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6622_ _6622_/A1 _6622_/A2 _6622_/B _7919_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_177_367 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_177_389 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6553_ hold90/Z _6553_/A2 _6553_/B _7901_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_3765_ _3765_/A1 _3765_/A2 _3765_/B _7973_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_173_551 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3696_ _7735_/Q _3696_/ZN VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_5504_ _5545_/A2 _5687_/B _5504_/A3 _5504_/B1 _5543_/B _5505_/A4 VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai32_1
X_6484_ hold469/Z _6485_/A2 _6485_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_145_286 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5435_ _5435_/A1 _5435_/A2 _5446_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_105_106 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
Xoutput310 _7941_/Q wb_ack_o VDD VSS gf180mcu_fd_sc_mcu7t5v0__buf_8
XFILLER_133_437 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xoutput332 _7947_/Q wb_dat_o[29] VDD VSS gf180mcu_fd_sc_mcu7t5v0__buf_8
Xoutput321 _7481_/Q wb_dat_o[19] VDD VSS gf180mcu_fd_sc_mcu7t5v0__buf_8
X_5366_ _4965_/B _5366_/A2 _4993_/C _5689_/A1 _5622_/A1 _5572_/C VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai32_1
X_5297_ _5006_/C _5709_/A2 _5297_/B _5378_/C _5299_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi211_1
X_4317_ _7414_/Q _4294_/Z _4317_/A3 _4318_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor3_1
XFILLER_141_492 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_7105_ _7105_/A1 _7105_/A2 _7105_/A3 _7105_/A4 _7106_/A4 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand4_1
XFILLER_59_215 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7036_ _7849_/Q _7193_/A2 _7189_/A2 _7711_/Q _7203_/B1 _7881_/Q _7039_/A2 VDD VSS
+ gf180mcu_fd_sc_mcu7t5v0__aoi222_1
X_4248_ _4248_/A1 _4248_/A2 _4248_/A3 _4248_/A4 _4283_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand4_2
XFILLER_142_37 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_68_771 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_28_602 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_67_292 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4179_ _4179_/A1 _4179_/A2 _4179_/A3 _4179_/A4 _4187_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand4_1
XFILLER_83_774 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_55_465 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1027 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1038 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_7938_ _7938_/D _7961_/RN _7938_/CLK _7938_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_43_638 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1005 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1016 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_150_6 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1049 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_148 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7869_ _7869_/D _7901_/RN _7877_/CLK _7869_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_23_373 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_168_389 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_149_570 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_137_721 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_167_56 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_109_456 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_164_584 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_152_702 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_137_776 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_3_712 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_152_757 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_151_212 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_78_502 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_4_2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_105_695 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_2_266 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_120_676 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_76_53 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_76_97 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_34_605 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2262 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2251 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2240 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_61_424 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_61_413 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2295 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2284 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2273 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
Xclkbuf_leaf_41_csclk clkbuf_3_7__f_csclk/Z _7743_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XTAP_1550 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_92_85 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_33_137 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1594 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1583 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1572 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1561 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_90 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
Xclkbuf_leaf_56_csclk clkbuf_3_6__f_csclk/Z _7819_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_127_242 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_143_702 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_5220_ _5538_/A1 _5042_/Z _5176_/B _5652_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_143_735 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_127_286 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5151_ _5151_/A1 _5151_/A2 _5024_/Z _5539_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_111_621 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_96_321 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_37_2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5082_ _5319_/C _5714_/B1 _5307_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_111_632 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_110_120 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4102_ _7808_/Q _6350_/A1 _4232_/A2 input5/Z _6418_/A1 _7840_/Q _4104_/A3 VDD VSS
+ gf180mcu_fd_sc_mcu7t5v0__aoi222_1
XFILLER_110_153 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4033_ _7664_/Q _6039_/A1 _4505_/A1 _7367_/Q _6333_/A1 _7802_/Q _4035_/A3 VDD VSS
+ gf180mcu_fd_sc_mcu7t5v0__aoi222_1
XFILLER_65_730 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_80_744 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_25_638 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5984_ hold278/Z _5987_/A2 _5985_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_7723_ _7723_/D _7901_/RN _7805_/CLK _7723_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
X_4935_ _5230_/A1 _5271_/A3 _5482_/B2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_2
XFILLER_21_811 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_178_676 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_138_507 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7654_ _7654_/D _7961_/RN _7694_/CLK _7654_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffsnq_1
XFILLER_20_321 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_4866_ hold668/Z _4867_/A2 _4867_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_177_197 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_177_175 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_138_529 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3817_ _3817_/I _4686_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_7585_ _7585_/D _7901_/RN _7691_/CLK _7585_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
X_4797_ _7230_/A1 _4795_/S _4797_/B _7485_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_6605_ _7914_/Q _7913_/Q _6950_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_4
X_6536_ hold90/Z _6536_/A2 _6536_/B _7893_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_21_26 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3748_ _7344_/Q _7411_/Q _3751_/A2 _3749_/S VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_180_318 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_137_26 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_119_776 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_133_212 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6467_ hold470/Z _6468_/A2 _6468_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_3679_ _7865_/Q _3679_/ZN VDD VSS gf180mcu_fd_sc_mcu7t5v0__inv_1
XFILLER_161_565 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5418_ _5692_/B _5563_/B2 _5618_/A3 _5419_/C VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor3_1
X_6398_ hold68/Z _6400_/A2 _6398_/B _7828_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_88_800 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xoutput195 _3681_/ZN mgmt_gpio_oeb[31] VDD VSS gf180mcu_fd_sc_mcu7t5v0__buf_8
X_5349_ _5482_/B2 _5510_/A2 _5493_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
Xoutput173 _3701_/ZN mgmt_gpio_oeb[11] VDD VSS gf180mcu_fd_sc_mcu7t5v0__buf_8
Xoutput184 _3691_/ZN mgmt_gpio_oeb[21] VDD VSS gf180mcu_fd_sc_mcu7t5v0__buf_8
XFILLER_0_737 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_102_632 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_87_354 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_102_676 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_101_153 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_7019_ _7880_/Q _7203_/B1 _7204_/A2 _7840_/Q _7832_/Q _7203_/A2 _7025_/A1 VDD VSS
+ gf180mcu_fd_sc_mcu7t5v0__aoi222_1
XFILLER_46_34 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_16_605 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_169_621 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_70_287 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_178_33 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_168_142 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_141_2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_51_490 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_62_99 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_11_354 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_137_540 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_164_392 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_109_286 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_127_70 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_11_70 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_140_738 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_608 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_619 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_78_321 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_19_421 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_93_357 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2070 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_62_766 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2092 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2081 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_99_4 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1391 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1380 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_4720_ hold724/Z _4731_/A2 _4721_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_4651_ _7457_/Q _3830_/Z _4651_/B _4652_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_175_657 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
Xinput31 mask_rev_in[5] input31/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
Xinput20 mask_rev_in[24] input20/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
Xinput64 mgmt_gpio_in[35] input64/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
Xinput42 mgmt_gpio_in[15] input42/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
Xinput53 mgmt_gpio_in[25] input53/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_7370_ _7370_/D _7961_/RN _7370_/CLK _7370_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffsnq_2
X_4582_ hold758/Z _4583_/A2 _4583_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
Xinput97 wb_adr_i[11] input97/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
X_6321_ hold137/Z _6332_/A2 hold138/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_115_223 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_115_212 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_115_201 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xinput86 spimemio_flash_io0_oeb input86/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_6_380 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xinput75 porb input75/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__buf_20
X_6252_ _4454_/Z _6264_/A2 _6252_/B _7759_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_5203_ _5203_/I _5375_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_6183_ hold73/Z _6191_/A2 _6183_/B _7727_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_5134_ _3723_/I _5777_/A1 _5538_/A1 _5026_/Z _5451_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__and4_1
XFILLER_97_641 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_69_321 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_69_354 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5065_ _5476_/B _5689_/A1 _5072_/B _5359_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_111_495 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_29_229 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_84_379 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4016_ _4013_/Z _4016_/A2 _4016_/A3 _4025_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_72_519 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_38_774 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_16_37 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5967_ hold347/Z _5970_/A2 _5968_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_52_276 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_53_799 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_4918_ _3722_/I _5006_/B _5006_/C _3728_/I _4945_/B1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand4_1
X_7706_ _7706_/D _7961_/RN _7706_/CLK _7706_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_21_630 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_178_495 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5898_ hold47/Z _5902_/A2 _5898_/B _7593_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_7637_ _7637_/D _7961_/RN _7643_/CLK _7637_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffsnq_1
XFILLER_20_140 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_21_641 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_166_646 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_138_337 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4849_ hold683/Z _4852_/A2 _4850_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_7568_ _7568_/D _7961_/RN _7587_/CLK _7568_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_181_638 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_146_392 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_134_521 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_106_212 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6519_ hold90/Z _6519_/A2 _6519_/B _7885_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_7499_ _7499_/D _7912_/CLK _7499_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_107_779 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_134_598 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_121_215 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_523 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_102_473 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_589 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_48_505 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_102_495 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_180_56 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_75_357 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_113_61 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_113_50 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_16_402 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_29_785 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_44_733 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_56_571 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_73_32 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_44_799 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_157_635 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_8_612 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_8_601 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_172_605 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_144_318 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_7_144 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_138_80 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_125_565 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_405 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_79_641 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_449 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_438 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_427 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_416 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_3_383 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_78_140 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_78_195 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_39_549 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_62_552 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_6870_ _7960_/Q _6880_/A2 _6893_/C1 _7472_/Q _6871_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_179_215 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5821_ _4454_/Z _5827_/A2 _5821_/B _7559_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_34_254 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5752_ _5777_/A1 _5608_/B _5752_/B1 _4996_/Z _5752_/C _5753_/C VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi221_1
XFILLER_50_747 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4703_ _7989_/I _4718_/A1 _4706_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_148_646 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_5683_ _5433_/C _5683_/A2 _5684_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_30_460 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4634_ _3830_/Z hold73/Z _4635_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_163_627 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_7422_ _7422_/D _7901_/RN _7849_/CLK _7996_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_163_649 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_162_137 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_162_115 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xhold612 _7384_/Q hold612/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
X_7353_ _7353_/D _7961_/RN _7353_/CLK _7353_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffsnq_2
Xhold601 hold601/I _7473_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
X_4565_ hold647/Z _4568_/A2 _4566_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
Xhold634 _7461_/Q hold634/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
XFILLER_128_392 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6304_ hold330/Z _6315_/A2 _6305_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
Xhold645 _7775_/Q hold645/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
Xhold623 hold623/I _7505_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
X_7284_ _7284_/I _7959_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_103_215 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
Xhold667 _7823_/Q hold667/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
X_4496_ hold73/Z _4504_/A2 _4496_/B hold557/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
Xhold678 _7387_/Q hold678/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
Xhold656 _7401_/Q hold656/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
X_6235_ hold302/Z _6242_/A2 _6236_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_134_16 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_131_546 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
Xhold689 _7677_/Q hold689/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
X_6166_ hold73/Z _6174_/A2 _6166_/B _7719_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_69_140 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_950 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_961 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_57_302 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5117_ _5392_/A1 _5344_/A2 _5680_/B2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_2
X_6097_ hold416/Z _6106_/A2 _6098_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_972 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_983 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_994 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_5048_ _5309_/A1 _3723_/I _5254_/A2 _5102_/B1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor3_1
XFILLER_84_132 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_57_357 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_150_37 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_84_187 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_84_176 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_25_210 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_26_744 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_13_405 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_25_254 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_53_563 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6999_ _7775_/Q _7200_/A2 _7201_/A2 _7749_/Q _7200_/B1 _7863_/Q _7000_/A4 VDD VSS
+ gf180mcu_fd_sc_mcu7t5v0__aoi222_1
XFILLER_138_101 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_166_421 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_159_79 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_154_605 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_138_156 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_126_318 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_147_690 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_181_457 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_104_2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_88_460 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_124_82 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_91_603 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_75_132 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_64_806 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_48_368 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_44_530 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_90_179 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_90_157 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_16_254 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_177_708 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_140_81 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_32_747 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_260 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_169_292 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_293 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_282 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_271 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_145_638 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_144_104 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_8_486 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_172_457 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4350_ _6567_/A1 _7905_/Q _6569_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_4_670 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_140_321 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_4281_ _4281_/A1 _4281_/A2 _4281_/A3 _4281_/A4 _4282_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor4_1
XFILLER_101_708 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6020_ hold336/Z _6021_/A2 _6021_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_140_387 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_67_622 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_94_463 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_39_357 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7971_ _7971_/D _7324_/Z _4415_/A2 _7971_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_66_176 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xclkbuf_3_3__f_csclk clkbuf_0_csclk/Z _7961_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
X_6922_ _6599_/Z _6955_/A4 _6908_/Z _7191_/B1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor3_4
XFILLER_81_168 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6853_ _7533_/Q _6878_/A2 _6853_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__or2_1
XFILLER_35_552 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_35_563 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5804_ _5804_/A1 _5804_/A2 _5804_/A3 _5804_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__or3_1
XFILLER_62_371 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_22_202 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_23_758 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_35_585 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6784_ _7649_/Q _6880_/C2 _6882_/A2 _7380_/Q _7819_/Q _6880_/A2 _6787_/A1 VDD VSS
+ gf180mcu_fd_sc_mcu7t5v0__aoi222_1
X_3996_ _3996_/A1 _3996_/A2 _3996_/A3 _3997_/C VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand3_1
X_5735_ _5104_/B _5735_/A2 _5247_/B _5724_/B _5735_/C _5736_/A4 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi221_2
XFILLER_31_780 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_50_599 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_176_763 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_136_605 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5666_ _5666_/A1 _5709_/A1 _5777_/A2 _5667_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_175_295 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_108_318 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7405_ _7405_/D _7961_/RN _7876_/CLK _7405_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
X_4617_ hold620/Z _4618_/A2 _4618_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_5597_ _5417_/I _5450_/C _5656_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_1
Xhold420 _7695_/Q hold420/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
X_4548_ hold90/Z _4548_/A2 _4548_/B _7382_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_144_682 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_144_671 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7336_ _7336_/D _7291_/Z _4031_/C2 _7336_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
Xhold442 _7656_/Q hold442/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
Xhold431 hold431/I _4482_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
Xhold453 _7352_/Q hold453/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
X_7267_ _7267_/A1 _7280_/A2 _7277_/B _7267_/C _7268_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi211_1
X_4479_ _7506_/Q _7273_/A1 hold67/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
Xhold464 _7828_/Q hold464/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
Xhold486 _7867_/Q hold486/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
Xhold475 _7877_/Q hold475/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
XFILLER_89_224 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6218_ hold487/Z _6225_/A2 _6219_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
Xhold497 _7650_/Q hold497/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
X_7198_ _7198_/A1 _7198_/A2 _7198_/A3 _7198_/A4 _7198_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__and4_1
X_6149_ hold73/Z _6157_/A2 _6149_/B _7711_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
XTAP_780 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_791 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_161_69 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_58_688 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_58_699 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_26_530 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1924 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1913 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1902 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_72_179 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1968 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1957 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1946 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1935 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_13_224 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_14_736 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_14_747 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1979 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_139_432 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_182_744 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_181_210 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_154_413 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_127_649 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_127_638 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_126_126 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_70_99 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_134_181 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_122_321 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_135_81 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_110_549 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_89_780 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_76_463 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_91_499 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_3850_ _3850_/A1 _3864_/A2 hold24/Z hold274/I hold133/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand4_4
XFILLER_158_741 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3781_ hold121/Z _7338_/Q _7414_/Q _3781_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_13_780 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_20_717 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_157_240 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_5520_ _5359_/B _5520_/A2 _5520_/B _5520_/C _5522_/B1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XFILLER_118_605 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_172_210 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_117_126 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_8_250 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5451_ _5774_/A1 _5643_/A2 _5451_/B _5460_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_67_2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5382_ _5022_/B _5205_/Z _5382_/A3 _5382_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__or3_1
XFILLER_114_811 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4402_ _4402_/A1 _4334_/Z _4402_/B _7334_/Q _4403_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XFILLER_141_641 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7121_ _7121_/A1 _7121_/A2 _7121_/A3 _7121_/A4 _7130_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand4_1
X_4333_ input67/Z _7582_/Q _4335_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_2
XFILLER_113_354 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7052_ _7647_/Q _7195_/A2 _7190_/B1 _7615_/Q _7053_/A4 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_4264_ _4264_/A1 _4264_/A2 _4264_/A3 _4264_/A4 _4281_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand4_1
XFILLER_115_29 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_113_398 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6003_ hold310/Z _6004_/A2 hold311/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_4195_ _7775_/Q _6282_/A1 _4888_/A1 _7536_/Q _6401_/A1 _7831_/Q _4198_/A2 VDD VSS
+ gf180mcu_fd_sc_mcu7t5v0__aoi222_1
XFILLER_95_783 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7954_ _7954_/D _7959_/RN _4411_/I1 hold39/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_131_39 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_55_636 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1209 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_6905_ _6905_/A1 _6905_/A2 _6941_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_4
XFILLER_54_179 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_7885_ _7885_/D _7901_/RN _7901_/CLK _7885_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_24_15 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6836_ _7821_/Q _6880_/A2 _6880_/B1 _7813_/Q _7651_/Q _6880_/C2 _6839_/A1 VDD VSS
+ gf180mcu_fd_sc_mcu7t5v0__aoi222_1
XFILLER_23_566 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_23_555 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_24_37 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_50_352 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6767_ _7736_/Q _6830_/B _6889_/A2 _7704_/Q _6767_/C _6771_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi221_1
XFILLER_10_205 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3979_ _7811_/Q _6350_/A1 _6333_/A1 _7803_/Q _3992_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_5718_ _5590_/B _5581_/B _5718_/A3 _5719_/A4 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor3_1
XFILLER_136_413 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_109_638 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6698_ _7637_/Q _6890_/A2 _6665_/Z _7741_/Q _6698_/C _6707_/B1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi221_1
XFILLER_164_744 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_163_232 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_136_457 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5649_ _5673_/A3 _5647_/B _5649_/A3 _5649_/A4 _5655_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand4_1
X_7319_ _7901_/RN _4334_/Z _7319_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__and2_1
Xhold250 hold250/I _7630_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
Xhold261 hold261/I _6254_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
XFILLER_117_682 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_104_321 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_6_6 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
Xhold283 _7729_/Q hold283/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
Xhold294 hold294/I _7663_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
Xhold272 _7343_/Q hold272/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
XFILLER_77_227 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_49_89 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_105_51 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_93_709 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_105_73 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_58_485 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_58_463 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2400 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_171_2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_45_113 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_73_466 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_65_77 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1743 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1732 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1721 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1710 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_73_499 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1776 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1765 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1754 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1798 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1787 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_155_700 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_127_424 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_182_585 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_170_769 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_170_747 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_135_490 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_107_181 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_5_286 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_30_91 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_123_641 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_1_492 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_77_783 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
Xinput7 mask_rev_in[12] input7/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_92_742 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_36_135 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_49_496 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_64_477 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4951_ _4951_/A1 _4951_/A2 _4951_/B _5016_/B _5602_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai211_4
XFILLER_17_382 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_36_179 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_177_302 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3902_ _7885_/Q _6503_/A1 _5903_/A1 input42/Z _4231_/B1 input70/Z _3906_/A1 VDD VSS
+ gf180mcu_fd_sc_mcu7t5v0__aoi222_1
X_7670_ _7670_/D _7961_/RN _7702_/CLK _7670_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffsnq_1
X_4882_ _4454_/Z _4882_/A2 _4882_/B _7532_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_177_313 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3833_ hold19/Z _3925_/A2 hold127/Z _3963_/A4 hold146/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand4_4
X_6621_ _7919_/Q _6621_/A2 _6622_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_177_357 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_146_700 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6552_ hold465/Z _6553_/A2 _6553_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_3764_ _3765_/A2 _3764_/A2 _3765_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_9_570 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3695_ _7743_/Q _3695_/ZN VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_5503_ _5797_/A2 _5546_/A2 _5546_/B1 _5543_/B _5503_/C _5509_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai221_1
XFILLER_146_744 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6483_ hold68/Z _6485_/A2 _6483_/B _7868_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_160_202 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5434_ _5789_/A1 _5614_/A3 _5625_/A2 _5434_/A4 _5435_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand4_1
Xoutput300 _4331_/Z serial_clock VDD VSS gf180mcu_fd_sc_mcu7t5v0__buf_8
XFILLER_105_118 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
Xoutput311 _7496_/Q wb_dat_o[0] VDD VSS gf180mcu_fd_sc_mcu7t5v0__buf_8
Xoutput322 _7497_/Q wb_dat_o[1] VDD VSS gf180mcu_fd_sc_mcu7t5v0__buf_8
Xoutput333 _7498_/Q wb_dat_o[2] VDD VSS gf180mcu_fd_sc_mcu7t5v0__buf_8
XFILLER_160_257 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5365_ _5797_/A1 _5099_/B _5365_/B1 _5681_/A1 _5408_/C VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai22_1
X_7104_ _7883_/Q _7203_/B1 _7204_/A2 _7843_/Q _7105_/A4 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_5296_ _5371_/C _5405_/B _5378_/C VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_4316_ _7337_/Q _7336_/Q _7338_/Q _4317_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_113_173 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_113_195 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_101_357 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7035_ _7035_/A1 _7035_/A2 _7035_/A3 _7035_/A4 _7035_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__and4_1
XFILLER_75_709 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4247_ _7676_/Q _6073_/A1 _5971_/A1 _7628_/Q _4248_/A4 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_4178_ _7759_/Q _6248_/A1 _4549_/A1 _7384_/Q _4179_/A4 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_95_580 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_67_282 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_27_146 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_28_669 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_70_414 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7937_ _7937_/D _7961_/RN _7938_/CLK _7937_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XTAP_1028 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_105 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_55_499 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_1006 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1017 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_7868_ _7868_/D _7901_/RN _7868_/CLK _7868_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XTAP_1039 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_6819_ _6819_/A1 _6819_/A2 _6819_/A3 _6819_/A4 _6825_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand4_1
XFILLER_51_672 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_156_519 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_156_508 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7799_ _7799_/D _7901_/RN _7799_/CLK _7799_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffsnq_1
XFILLER_51_24 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_51_57 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_167_68 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_152_747 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_124_438 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_151_246 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_105_641 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_3_779 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_3_757 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_116_50 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_105_685 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_104_162 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_59_783 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_19_636 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2252 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2241 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2230 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_92_53 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_18_179 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2296 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2285 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2274 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2263 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_159_302 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1551 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1540 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_61_458 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1584 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1573 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1562 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_30_812 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_80 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_91 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_159_357 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1595 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_128_744 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_128_755 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_127_210 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_182_360 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_6_540 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_115_438 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_130_408 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_170_599 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5150_ _5151_/A1 _5151_/A2 _5024_/Z _5150_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__and3_1
XFILLER_151_780 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_97_812 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5081_ _4898_/Z _5254_/A3 _5714_/B1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_2
XFILLER_110_132 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4101_ input37/Z _5903_/A1 _4488_/A1 _7357_/Q _5874_/A1 _7583_/Q _4104_/A2 VDD VSS
+ gf180mcu_fd_sc_mcu7t5v0__aoi222_1
XFILLER_96_333 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_57_709 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_111_699 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_110_165 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_4032_ _4032_/A1 _4032_/A2 _4036_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_77_580 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_65_720 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5983_ hold47/Z _5987_/A2 _5983_/B hold282/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_65_797 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_24_105 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_24_116 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_37_499 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_178_600 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4934_ _5199_/B _5201_/B _5271_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_4
X_7722_ _7722_/D _7901_/RN _7820_/CLK _7722_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_177_110 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_166_806 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4865_ _4448_/Z _4867_/A2 _4865_/B _7525_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_7653_ _7653_/D _7961_/RN _7733_/CLK _7653_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffsnq_1
X_3816_ hold123/Z _3925_/A2 hold127/Z _3794_/Z _3817_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__or4_4
X_7584_ _7584_/D _7901_/RN _7691_/CLK _7584_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
X_4796_ _7485_/Q _4795_/S _4797_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_6604_ _7913_/Q _6609_/A2 _6604_/B _7913_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_6535_ hold466/Z _6536_/A2 _6536_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_3747_ _4284_/A1 _3763_/B _3747_/B _7977_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_20_399 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_137_16 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_161_511 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_134_747 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_118_276 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3678_ _7873_/Q _3678_/ZN VDD VSS gf180mcu_fd_sc_mcu7t5v0__inv_1
XFILLER_106_449 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_106_438 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_106_427 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6466_ hold68/Z _6468_/A2 _6466_/B _7860_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_5417_ _5417_/I _5446_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_6397_ hold464/Z _6400_/A2 _6398_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
Xoutput174 _3700_/ZN mgmt_gpio_oeb[12] VDD VSS gf180mcu_fd_sc_mcu7t5v0__buf_8
Xoutput185 _3690_/ZN mgmt_gpio_oeb[22] VDD VSS gf180mcu_fd_sc_mcu7t5v0__buf_8
X_5348_ _5685_/B _5624_/A2 _5642_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
Xoutput196 _3680_/ZN mgmt_gpio_oeb[32] VDD VSS gf180mcu_fd_sc_mcu7t5v0__buf_8
X_7018_ _7750_/Q _7201_/A2 _7201_/B1 _7670_/Q _7023_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_5279_ _5616_/A1 _5237_/Z _5712_/B _5573_/B _5282_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XFILLER_83_583 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_71_712 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_43_425 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_102_52 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_62_34 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_12_812 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_30_108 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_178_56 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_168_176 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_134_2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_7_304 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_23_193 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_7_359 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_125_736 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_124_213 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_127_60 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_3_554 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_152_599 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_105_460 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_79_812 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_3_587 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_609 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_87_75 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_39_709 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_120_463 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_93_303 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_19_499 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_2060 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2093 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2082 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2071 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1392 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1381 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1370 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_30_620 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_147_327 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4650_ _3830_/Z hold90/Z _4651_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_1
Xinput10 mask_rev_in[15] input10/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
Xinput21 mask_rev_in[25] input21/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_174_179 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xinput43 mgmt_gpio_in[16] input43/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
Xinput54 mgmt_gpio_in[26] input54/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_6320_ _4454_/Z _6332_/A2 _6320_/B _7791_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
Xinput32 mask_rev_in[6] input32/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_4581_ _4448_/Z _4583_/A2 _4581_/B _7395_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
Xinput98 wb_adr_i[12] input98/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
Xinput65 mgmt_gpio_in[36] _8008_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_128_585 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_116_747 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xinput87 spimemio_flash_io1_do _8007_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
Xinput76 qspi_enabled _4387_/S VDD VSS gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_143_566 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_115_246 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6251_ hold644/Z _6264_/A2 _6252_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_6_392 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5202_ _5202_/A1 _5202_/A2 _5371_/B _5371_/C _5203_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_2
X_6182_ hold331/Z _6191_/A2 _6183_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_88_108 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5133_ _5309_/A1 _3723_/I _5394_/A1 _5006_/C _5645_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand4_4
XFILLER_69_344 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_69_377 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5064_ _5301_/A1 _5062_/Z _5064_/B _5072_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_96_174 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_57_539 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4015_ _7672_/Q _6056_/A1 _5886_/A1 input56/Z _5817_/A1 _7562_/Q _4016_/A3 VDD VSS
+ gf180mcu_fd_sc_mcu7t5v0__aoi222_1
XFILLER_25_425 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_53_712 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_80_531 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_37_296 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_12_108 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_5966_ hold47/Z _5970_/A2 _5966_/B hold360/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_52_266 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4917_ _3722_/I _5006_/B _5006_/C _3728_/I _4917_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__and4_2
X_7705_ _7705_/D _7961_/RN _7735_/CLK _7705_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
X_5897_ hold526/Z _5902_/A2 _5898_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_178_463 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7636_ _7636_/D _7961_/RN _7643_/CLK _7636_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffsnq_1
X_4848_ _4848_/A1 _7285_/A2 _4852_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_32_37 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_165_113 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_148_37 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_21_697 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_180_105 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_107_703 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4779_ _4779_/A1 _7285_/A2 _4783_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_7567_ _7567_/D input75/Z _7567_/CLK _7567_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffsnq_2
XFILLER_107_725 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6518_ hold462/Z _6519_/A2 _6519_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_4_318 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7498_ _7498_/D _7912_/CLK _7498_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_6449_ hold68/Z _6451_/A2 _6449_/B hold290/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
Xclkbuf_leaf_40_csclk clkbuf_3_7__f_csclk/Z _7816_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_102_463 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_102_441 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_87_141 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_48_517 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_102_485 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_57_67 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xclkbuf_leaf_55_csclk clkbuf_3_6__f_csclk/Z _7698_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_57_89 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_113_73 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_16_458 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_44_756 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_31_428 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_11_141 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_169_496 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_12_686 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_22_70 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_156_179 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_152_330 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_180_672 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_152_385 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_113_728 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_406 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_79_620 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_439 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_428 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_417 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_79_653 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_121_783 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_93_144 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_93_155 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_93_177 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_35_712 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_62_542 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_62_531 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_62_564 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5820_ hold626/Z _5827_/A2 _5821_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_50_704 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5751_ _5778_/A1 _5776_/A3 _5776_/A4 _5754_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_97_2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_50_759 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4702_ _4718_/A1 hold168/Z _4702_/B hold169/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_7421_ hold62/Z _7901_/RN _7816_/CLK _7995_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_147_135 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5682_ _5682_/A1 _5692_/A2 _5682_/A3 _5683_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand3_1
X_4633_ _7993_/I _4652_/A1 _4636_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_147_146 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_175_499 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_118_29 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_116_500 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7352_ _7352_/D _7961_/RN _7353_/CLK _7352_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffsnq_1
Xhold602 _7510_/Q hold602/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
X_4564_ _4564_/A1 _7285_/A2 _4568_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_7283_ hold31/I _7517_/Q _7279_/B _7283_/B _7284_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai31_1
Xmax_cap343 hold32/Z _7285_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__buf_20
X_6303_ _4454_/Z _6315_/A2 _6303_/B _7783_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
Xhold624 _7692_/Q hold624/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
Xhold635 _7445_/Q hold635/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
Xhold613 _7398_/Q hold613/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
X_6234_ hold73/Z _6242_/A2 _6234_/B _7751_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_131_503 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_89_428 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xhold646 _7783_/Q hold646/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
Xhold679 _7468_/Q hold679/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
X_4495_ hold555/Z _4504_/A2 hold556/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
Xhold668 _7526_/Q hold668/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
Xhold657 _7831_/Q hold657/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
X_6165_ hold333/Z _6174_/A2 _6166_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_134_28 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_97_461 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_85_601 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_940 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_951 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_962 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_5116_ _5309_/A1 _3723_/I _5344_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_2
XFILLER_97_494 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6096_ _4460_/Z _6106_/A2 _6096_/B _7686_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_85_645 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_973 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_984 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_995 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_5047_ _5006_/B _5254_/A2 _5254_/A3 _5689_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand3_4
XFILLER_45_509 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_27_48 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_150_49 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_53_531 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_6998_ _7823_/Q _7202_/A2 _7202_/B1 _7783_/Q _7759_/Q _7202_/C2 _7000_/A3 VDD VSS
+ gf180mcu_fd_sc_mcu7t5v0__aoi222_1
X_5949_ hold47/Z _5953_/A2 _5949_/B hold429/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_13_439 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_13_428 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_179_783 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_40_247 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_159_69 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7619_ _7619_/D _7961_/RN _7698_/CLK _7619_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_181_425 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_175_13 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_138_179 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_5_638 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_161_160 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_150_812 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_68_33 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_321 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_130_580 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_103_783 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_88_494 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_76_623 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_387 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_124_50 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_102_282 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_75_144 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_90_103 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_84_54 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_75_177 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_75_155 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_17_712 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_17_70 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_169_260 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_261 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_250 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_90_9 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_31_247 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_294 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_283 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_272 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_12_450 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_172_414 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_157_499 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_172_469 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_137_190 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_99_704 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_141_812 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_140_333 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_98_247 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4280_ _4280_/A1 _4280_/A2 _4274_/Z _4279_/Z _4281_/A4 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand4_1
XFILLER_121_580 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_79_494 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_79_483 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_66_100 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_39_303 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_12_2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7970_ _7970_/D _7323_/Z _4415_/A2 _7970_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_94_475 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_66_166 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_54_317 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6921_ _7660_/Q _7194_/B1 _6959_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_66_188 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6852_ _7133_/S _6852_/A2 _6852_/B _7928_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_5803_ _5803_/A1 _5803_/A2 _5803_/A3 _5803_/A4 _5804_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand4_1
XFILLER_50_534 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6783_ _6879_/A1 _6783_/A2 _6793_/C VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_3995_ _7859_/Q _6452_/A1 _5988_/A1 _7641_/Q _3995_/C _3999_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi221_4
XFILLER_22_247 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_50_556 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_5734_ _5778_/A1 _5733_/Z _5737_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_5665_ _5665_/A1 _5753_/B _5671_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_163_425 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7404_ _7404_/D _7961_/RN _7874_/CLK _7404_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
X_4616_ _4448_/Z _4618_/A2 _4616_/B _7409_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_5596_ _5448_/B _5596_/A2 _5661_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_1
Xhold410 _7781_/Q hold410/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
X_7335_ _7335_/D _7290_/Z _4418_/I1 _7335_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
X_4547_ hold217/Z _4548_/A2 _4548_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_150_108 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_132_812 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xhold421 _7819_/Q hold421/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
Xhold443 hold443/I _7656_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
Xhold432 hold432/I _7353_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
Xhold454 hold454/I _4477_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
X_7266_ _7266_/A1 _7266_/A2 _7267_/C VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
Xhold487 _7744_/Q hold487/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
XFILLER_143_193 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xhold465 _7901_/Q hold465/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
Xhold476 _7359_/Q hold476/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
X_4478_ hold430/Z _4487_/A1 hold431/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_6217_ hold73/Z _6225_/A2 _6217_/B _7743_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
Xhold498 hold498/I _7650_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
X_7197_ _7536_/Q _7197_/A2 _6938_/I _7392_/Q _7198_/A4 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_6148_ hold307/Z _6157_/A2 _6149_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_770 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_781 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_792 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_57_144 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_6079_ _4460_/Z _6089_/A2 _6079_/B hold216/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_85_464 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1925 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1914 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1903 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_159_709 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_159_4 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1958 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1947 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1936 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_41_534 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_54_68 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_1969 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_80_191 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_179_580 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_179_591 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_110_63 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_70_34 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_139_499 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_126_105 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_119_61 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_135_650 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_123_812 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_119_94 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_1_641 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_122_399 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_95_20 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_49_623 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_95_64 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_95_53 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_64_615 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_76_497 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_64_659 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_72_670 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_17_586 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_177_528 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_149_208 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_32_534 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3780_ _4291_/B _3780_/A2 _7962_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_173_712 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_145_425 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5450_ _5643_/A2 _5608_/B _5752_/B1 _4996_/Z _5450_/C _5461_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi221_1
XFILLER_117_116 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_9_785 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4401_ _7425_/Q _4334_/Z _4402_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_5381_ _5022_/B _5381_/A2 _5382_/A3 _5381_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__or3_1
XFILLER_173_778 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_145_469 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_132_108 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_126_672 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_153_491 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_141_631 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_125_171 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7120_ _7860_/Q _6938_/I _7188_/A2 _7381_/Q _7121_/A4 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_4332_ _4292_/B _3738_/Z _4291_/B _4382_/A2 _7411_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai22_1
XFILLER_5_73 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_99_567 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_87_707 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7051_ _7793_/Q _7190_/A2 _7190_/C1 _7703_/Q _7053_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_4263_ _4263_/A1 _4263_/A2 _4263_/A3 _4263_/A4 _4282_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor4_1
XFILLER_140_174 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_140_152 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6002_ hold68/Z _6004_/A2 _6002_/B hold341/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_67_442 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_28_807 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4194_ _4194_/A1 _4194_/A2 _4194_/A3 _4194_/A4 _4202_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand4_1
XFILLER_94_250 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_39_144 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_7953_ _7953_/D _7959_/RN _4411_/I1 hold71/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
X_6904_ _6955_/A4 _6941_/A1 _7202_/C2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_4
XFILLER_54_169 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_7884_ _7884_/D _7901_/RN _7900_/CLK _7884_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
X_6835_ _7643_/Q _6890_/A2 _6665_/Z _7747_/Q _6835_/C _6849_/B1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi221_1
XFILLER_50_331 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_149_720 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_6766_ _6766_/A1 _6766_/A2 _6766_/A3 _6766_/A4 _6777_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand4_1
X_3978_ _7875_/Q _6486_/A1 _5828_/A1 _7568_/Q _3994_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_50_364 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5717_ _5717_/A1 _5717_/A2 _5717_/A3 _5718_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor3_1
XFILLER_108_105 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xclkbuf_2_1__f_mgmt_gpio_in[4] clkbuf_0_mgmt_gpio_in[4]/Z _7977_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
X_6697_ _6697_/A1 _6697_/A2 _6697_/A3 _6698_/C VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_164_756 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5648_ _5648_/A1 _5648_/A2 _5624_/B _5648_/B2 _5648_/C _5743_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi221_1
XFILLER_40_37 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_156_37 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5579_ _5669_/A1 _5027_/Z _5579_/B _5710_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_105_812 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xhold251 _7754_/Q hold251/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
Xhold240 _7812_/Q hold240/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
XFILLER_151_428 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xhold262 hold262/I _7760_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
X_7318_ input75/Z _4334_/Z _7318_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__and2_1
X_7249_ _7519_/Q _7249_/A2 _7251_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
Xhold284 _7713_/Q hold284/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
Xhold295 _7665_/Q hold295/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
Xhold273 _3812_/Z hold273/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
XFILLER_131_141 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_77_239 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2401 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_45_125 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1700 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_164_2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1733 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1722 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1711 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_121_62 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_73_489 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_1766 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1755 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1744 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_121_73 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_81_33 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_14_534 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1799 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1777 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1788 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_41_353 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_41_397 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_167_561 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_155_712 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_182_542 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_154_211 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_10_784 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_6_744 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_5_221 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_154_266 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_114_108 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_182_597 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_135_480 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_107_160 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_110_325 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_1_482 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_76_250 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xinput8 mask_rev_in[13] input8/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_49_453 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_49_475 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_37_637 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_91_231 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4950_ _5069_/A2 _4930_/Z _5458_/C _5015_/B _5357_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XFILLER_91_286 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_17_361 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_51_106 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3901_ _3901_/A1 _3901_/A2 _3901_/A3 _3901_/A4 _3917_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand4_1
X_4881_ hold606/Z _4882_/A2 _4882_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_3832_ hold275/Z _3886_/A2 _6520_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_4
X_6620_ _7001_/C _4331_/Z _6621_/A2 _6620_/B _7918_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai31_1
XFILLER_32_353 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6551_ hold68/Z _6553_/A2 _6551_/B _7900_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_158_583 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5502_ _5502_/A1 _5652_/A3 _5767_/A2 _5641_/A2 _5509_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand4_1
X_3763_ _7973_/Q _7411_/Q _3763_/B _3764_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_3694_ _7751_/Q _3694_/ZN VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_6482_ hold458/Z _6485_/A2 _6483_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_5433_ _5062_/Z _5176_/B _5624_/B _5482_/B2 _5433_/C _5434_/A4 VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai221_1
Xoutput301 _3961_/Z serial_data_1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__buf_8
XFILLER_161_737 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_133_428 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_126_480 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5364_ _5669_/A1 _5608_/B _5573_/A1 _5292_/B _5732_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_1
Xoutput334 _7948_/Q wb_dat_o[30] VDD VSS gf180mcu_fd_sc_mcu7t5v0__buf_8
Xoutput323 _7482_/Q wb_dat_o[20] VDD VSS gf180mcu_fd_sc_mcu7t5v0__buf_8
Xoutput312 _7488_/Q wb_dat_o[10] VDD VSS gf180mcu_fd_sc_mcu7t5v0__buf_8
XFILLER_160_247 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4315_ _7338_/Q _4309_/S _4319_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_7103_ _7835_/Q _7203_/A2 _7204_/B1 _7771_/Q _7105_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_5295_ _5392_/A1 _5392_/A2 _5376_/B _5297_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor3_1
XFILLER_113_141 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_113_185 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_101_347 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7034_ _7751_/Q _7201_/A2 _7196_/A2 _7889_/Q _7035_/A4 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_4246_ _7814_/Q hold134/I _7285_/A1 _7960_/Q _4248_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_95_570 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_4177_ _7372_/Q _4522_/A1 _4574_/A1 _7394_/Q _7404_/Q _4599_/A1 _4179_/A3 VDD VSS
+ gf180mcu_fd_sc_mcu7t5v0__aoi222_1
XFILLER_83_732 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_55_412 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_55_445 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_7936_ _7936_/D _7961_/RN _7949_/CLK _7936_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XTAP_1029 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1018 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_43_629 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1007 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_169_804 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7867_ _7867_/D _7901_/RN _7867_/CLK _7867_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_168_325 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_168_303 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6818_ _7820_/Q _6880_/A2 _6893_/C1 _7634_/Q _6819_/A4 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_7798_ _7798_/D _7901_/RN _7802_/CLK _7798_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffsnq_1
XFILLER_137_712 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6749_ _7801_/Q _6883_/A2 _6883_/B1 _7785_/Q _6752_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_51_69 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_164_531 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_164_542 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_109_425 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_137_767 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_136_266 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_151_225 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_105_697 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_104_152 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_116_62 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_76_33 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_120_667 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_58_250 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_46_423 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_18_136 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2253 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2242 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2231 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2220 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_73_286 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2286 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2275 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2264 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1541 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1530 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2297 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1585 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1574 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1563 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1552 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_70 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_81 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_42_673 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_92 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_1596 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_14_386 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_6_530 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_170_534 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_115_428 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_51_6 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_142_247 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_108_491 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5080_ _5392_/A1 _5005_/Z _5779_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_2
X_4100_ _4100_/A1 _4100_/A2 _4100_/A3 _4100_/A4 _4105_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand4_1
XFILLER_84_518 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_4031_ _7786_/Q _6299_/A1 _4444_/A1 _7351_/Q _4231_/B1 _4031_/C2 _4032_/A2 VDD VSS
+ gf180mcu_fd_sc_mcu7t5v0__aoi222_1
XFILLER_77_592 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_77_570 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_49_283 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_37_467 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5982_ hold281/Z _5987_/A2 _5983_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_37_478 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_52_415 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4933_ _4917_/Z _4919_/Z _5201_/B _4941_/C VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi21_4
X_7721_ _7721_/D _7901_/RN _7819_/CLK _7721_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_24_139 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_52_459 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_177_144 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4864_ hold749/Z _4867_/A2 _4865_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_7652_ _7652_/D _7961_/RN _7733_/CLK _7652_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffsnq_1
X_7583_ hold33/Z _7901_/RN _7583_/CLK _7583_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_119_712 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_119_701 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3815_ _3796_/Z hold275/Z _6503_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_4
X_4795_ _7228_/I0 _7484_/Q _4795_/S _7484_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_20_345 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_32_194 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_6603_ _7913_/Q _6586_/B _6609_/A2 _6604_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_158_380 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_146_520 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_118_211 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6534_ hold68/Z _6536_/A2 _6534_/B _7892_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_3746_ input58/Z _7411_/Q _3763_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_20_389 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_180_309 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6465_ hold509/Z _6468_/A2 _6466_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_173_372 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5416_ _3722_/I _5709_/A1 _5452_/C _5543_/C _5417_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor4_4
X_3677_ _7932_/Q _7003_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_161_567 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_134_759 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6396_ hold47/Z _6400_/A2 _6396_/B _7827_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_5347_ _5768_/A2 _5680_/B1 _5347_/B _5347_/C _5353_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi211_1
Xoutput175 _3699_/ZN mgmt_gpio_oeb[13] VDD VSS gf180mcu_fd_sc_mcu7t5v0__buf_8
Xoutput186 _3689_/ZN mgmt_gpio_oeb[23] VDD VSS gf180mcu_fd_sc_mcu7t5v0__buf_8
XFILLER_0_717 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
Xoutput197 _3679_/ZN mgmt_gpio_oeb[33] VDD VSS gf180mcu_fd_sc_mcu7t5v0__buf_8
XFILLER_99_183 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5278_ _5292_/B _5724_/B _5363_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_7017_ _7776_/Q _7200_/A2 _7200_/B1 _7864_/Q _7023_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_101_144 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4229_ _7527_/Q _4868_/A1 _4893_/A1 _7537_/Q _4236_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_28_467 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_43_404 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_46_69 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_55_286 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_70_245 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7919_ _7919_/D _7961_/RN _7940_/CLK _7919_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_24_673 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_156_328 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_127_2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_109_233 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_180_810 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_152_534 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_124_247 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_3_544 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_140_729 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_87_21 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_133_792 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_59_570 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_47_721 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_62_713 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_2061 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2050 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_61_212 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2094 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2083 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2072 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_159_144 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1393 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1382 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1360 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1371 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_174_103 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_128_531 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xinput11 mask_rev_in[16] input11/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
Xinput22 mask_rev_in[26] input22/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_4580_ hold669/Z _4583_/A2 _4581_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_30_676 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_162_309 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
Xinput44 mgmt_gpio_in[17] input44/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
Xinput55 mgmt_gpio_in[27] input55/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
Xinput33 mask_rev_in[7] input33/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
Xinput66 mgmt_gpio_in[37] _8009_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_128_575 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
Xinput88 spimemio_flash_io1_oeb input88/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
Xinput77 ser_tx input77/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
Xinput99 wb_adr_i[13] input99/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
X_6250_ _4448_/Z _6264_/A2 _6250_/B _7758_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_5201_ _5200_/B _5230_/A1 _5663_/A1 _5201_/B _5371_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai31_1
XFILLER_170_353 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6181_ _4460_/Z _6191_/A2 _6181_/B hold120/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_42_2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5132_ _3722_/I _5087_/C _5006_/B _5254_/A2 _5643_/B1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor4_4
XFILLER_96_142 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5063_ _5006_/C _5616_/A1 _5563_/B2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_4
XFILLER_97_698 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_96_164 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_57_529 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_4014_ input30/Z _4249_/A2 _4232_/A2 input7/Z _6401_/A1 _7834_/Q _4016_/A2 VDD VSS
+ gf180mcu_fd_sc_mcu7t5v0__aoi222_1
XFILLER_25_415 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_92_392 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_25_448 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_37_286 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5965_ hold359/Z _5970_/A2 _5966_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_4916_ _3728_/I _5369_/B _5230_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_4
X_5896_ hold41/Z _5902_/A2 _5896_/B _7592_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_7704_ _7704_/D _7961_/RN _7704_/CLK _7704_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_21_621 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7635_ _7635_/D _7901_/RN _7806_/CLK _7635_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
X_4847_ _4454_/Z _4847_/A2 _4847_/B hold583/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_181_618 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_120_9 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_5_809 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4778_ _4454_/Z _4778_/A2 _4778_/B hold593/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_7566_ _7566_/D input75/Z _7567_/CLK _7566_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_180_128 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3729_ _5369_/B _5022_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_8
XFILLER_174_692 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_6517_ hold68/Z _6519_/A2 _6517_/B _7884_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_7497_ _7497_/D _7912_/CLK _7497_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_6448_ hold289/Z _6451_/A2 _6449_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_134_534 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_106_247 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_164_37 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_122_729 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6379_ hold47/Z _6383_/A2 _6379_/B _7819_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_102_431 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_88_676 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_87_153 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_558 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_102_475 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_180_58 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_75_348 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_90_318 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_83_392 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_71_565 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_43_256 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_12_676 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_22_60 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_171_128 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_165_692 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_138_93 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_152_375 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_125_567 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_429 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_418 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_407 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_94_602 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_120_250 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_78_197 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_19_242 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_74_392 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_62_521 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_19_286 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_62_576 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_35_779 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_179_239 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5750_ _5754_/A1 _5754_/A2 _5775_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_4701_ hold167/Z _3819_/Z _4701_/B hold168/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_5681_ _5681_/A1 _5620_/B _5681_/B _5723_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
XTAP_1190 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_175_423 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4632_ _4652_/A1 hold95/Z _4632_/B hold96/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_7420_ hold65/Z _7901_/RN _7816_/CLK _7994_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_30_451 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_175_456 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_162_128 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_156_670 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_7351_ _7351_/D _7961_/RN _7570_/CLK _7351_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffsnq_2
X_4563_ _4454_/Z _4563_/A2 _4563_/B _7388_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
Xhold603 hold603/I _7510_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
X_7282_ _7282_/A1 _7282_/A2 _7282_/B _7283_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_143_342 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_116_534 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xhold625 _7684_/Q hold625/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
X_6302_ hold646/Z _6315_/A2 _6303_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_4494_ _4460_/Z _4504_/A2 _4494_/B hold229/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
Xhold636 _7645_/Q hold636/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
Xhold614 _7372_/Q hold614/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
X_6233_ hold303/Z _6242_/A2 _6234_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
Xhold658 _7537_/Q hold658/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
Xhold669 _7395_/Q hold669/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
Xhold647 _7389_/Q hold647/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
XFILLER_170_183 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_143_386 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6164_ _4460_/Z _6174_/A2 _6164_/B hold147/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
XTAP_930 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_941 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_952 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_5115_ _4999_/Z _5115_/A2 _5474_/B _5361_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_6095_ hold199/Z _6106_/A2 _6096_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_963 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_974 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_985 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_996 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_5046_ _5709_/A1 _5005_/Z _5404_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_111_294 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_111_283 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_57_337 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_72_329 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_72_318 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_38_573 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_84_189 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_65_392 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_25_212 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_13_407 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_25_256 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6997_ _6997_/A1 _6997_/A2 _6997_/A3 _6997_/A4 _6997_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__and4_1
X_5948_ hold428/Z _5953_/A2 _5949_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_178_250 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_166_401 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_159_37 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_138_125 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5879_ hold653/Z _5880_/A2 _5880_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_7618_ _7618_/D _7961_/RN _7698_/CLK _7618_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_4_105 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7549_ _7549_/D _7308_/Z _4418_/I1 _7549_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffnrnq_1
XFILLER_175_47 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_146_191 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_119_383 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_162_673 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_122_515 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_107_567 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_161_172 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_122_526 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_1_812 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_68_56 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_49_805 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_102_250 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_75_112 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_124_62 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_17_702 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_91_638 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_56_370 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_56_392 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_71_351 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_31_215 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_251 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_240 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_169_283 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_295 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_284 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_273 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_262 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_129_125 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_33_70 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_157_456 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_149_70 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_8_433 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_138_692 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_125_353 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_4_661 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_180_481 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_79_451 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_79_440 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_140_389 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_121_570 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_121_592 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_82_605 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_82_638 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6920_ _6953_/A1 _6953_/A2 _6941_/A2 _7194_/B1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor3_4
XFILLER_23_705 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6851_ _7928_/Q _7133_/S _6852_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_5802_ _5802_/A1 _5802_/A2 _5806_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_6782_ _7737_/Q _6878_/A2 _6783_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_3994_ _3994_/A1 _3994_/A2 _3994_/A3 _3995_/C VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand3_2
XFILLER_16_790 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_50_546 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5733_ _5733_/A1 _5733_/A2 _5733_/A3 _5733_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__and3_1
XFILLER_148_445 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_129_29 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5664_ _5752_/B1 _5774_/A2 _5774_/B1 _5774_/A1 _5753_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_175_286 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5595_ _5661_/A1 _5662_/A1 _5319_/C _5596_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor3_1
XFILLER_135_117 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xclkbuf_leaf_54_csclk clkbuf_3_6__f_csclk/Z _7707_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
X_7403_ _7403_/D _7961_/RN _7871_/CLK _7403_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
X_4615_ hold711/Z _4618_/A2 _4616_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_4546_ hold68/Z _4548_/A2 _4546_/B _7381_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
Xhold411 _7826_/Q hold411/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
Xhold400 hold400/I _7370_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
X_7334_ _7334_/D _4440_/Z _7977_/CLK _7334_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_144_673 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_144_651 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
Xhold444 _7818_/Q hold444/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
Xhold422 _7721_/Q hold422/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
Xhold433 _7697_/Q hold433/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
X_7265_ _7518_/Q _7265_/A2 _7265_/B1 _7519_/Q _7266_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_116_375 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xhold466 _7893_/Q hold466/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
XFILLER_89_226 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_89_215 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xhold477 hold477/I _4498_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
X_4477_ _4487_/A1 hold47/Z _4477_/B hold455/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
Xhold455 hold455/I _7352_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
X_6216_ hold328/Z _6225_/A2 _6217_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
Xhold499 _7762_/Q hold499/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
Xclkbuf_leaf_69_csclk _7961_/CLK _7649_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
Xhold488 _7566_/Q hold488/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
X_7196_ _7547_/Q _7196_/A2 _7196_/B1 _7475_/Q _7198_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_6147_ _4460_/Z _6157_/A2 _6147_/B hold129/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_58_602 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_760 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_57_101 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_161_38 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_97_292 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_58_657 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_771 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_782 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_38_37 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_793 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_6078_ hold215/Z _6089_/A2 _6079_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_57_156 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5029_ _5643_/A2 _5027_/Z _5585_/B _5038_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_73_638 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_72_104 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1915 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1904 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_38_392 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1959 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1948 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1937 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1926 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_13_215 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_14_738 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_179_570 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_110_86 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_110_75 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_182_702 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_22_782 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_154_415 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_21_292 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_182_768 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_181_212 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_5_425 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_182_779 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_119_73 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_5_469 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_122_323 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_1_620 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_150_676 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_122_389 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_103_570 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_95_43 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_174 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_64_605 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_48_167 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_29_370 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_17_565 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_72_660 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_60_800 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_17_576 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_44_80 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_9_720 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_158_765 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_157_231 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_12_270 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_172_212 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_157_286 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_4400_ _7430_/Q input77/Z _4400_/S _4400_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_5380_ _5380_/I _5641_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_114_802 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_5_30 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_125_183 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_99_513 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4331_ _7918_/Q _7575_/Q _7580_/Q _4331_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_141_643 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_140_120 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_7050_ _7841_/Q _7204_/A2 _7204_/B1 _7769_/Q _7053_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_4262_ _4262_/A1 _4262_/A2 _4262_/A3 _4262_/A4 _4263_/A4 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand4_1
XFILLER_140_164 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6001_ hold340/Z _6004_/A2 _6002_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_79_281 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_67_432 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4193_ input53/Z _5886_/A1 _4759_/A1 _7469_/Q _4194_/A4 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_95_785 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_67_465 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_67_476 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_39_156 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7952_ _7952_/D _7959_/RN _4411_/I1 hold28/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_67_487 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_48_690 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_54_104 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_55_638 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6903_ _6908_/A1 _7913_/Q _6936_/A1 _6941_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand3_4
X_7883_ _7883_/D _7901_/RN _7883_/CLK _7883_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
X_6834_ _6834_/A1 _6834_/A2 _6834_/A3 _6834_/A4 _6835_/C VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand4_1
XFILLER_50_321 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_50_343 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6765_ _7752_/Q _6644_/Z _6665_/Z _7744_/Q _6891_/C1 _7778_/Q _6766_/A4 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi222_1
X_3977_ _7787_/Q _6299_/A1 _4219_/A2 input17/Z _3994_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_50_354 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5716_ _5716_/A1 _5716_/A2 _5716_/A3 _5732_/A3 _5717_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand4_1
XFILLER_50_387 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6696_ _7847_/Q _6890_/B1 _6894_/C1 _7831_/Q _6697_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_163_212 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5647_ _4993_/B _5647_/A2 _5741_/A3 _5647_/B _5648_/C VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai31_1
X_5578_ _5578_/A1 _5578_/A2 _5578_/A3 _5578_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__and3_1
Xhold252 _7730_/Q hold252/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
Xhold230 _7813_/Q hold230/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
Xhold241 _7560_/Q hold241/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
X_7317_ input75/Z _4334_/Z _7317_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__and2_1
X_4529_ _4448_/Z _4531_/A2 _4529_/B _7373_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_7248_ _7248_/A1 _7277_/B _7248_/B _7951_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi21_1
Xhold285 _7753_/Q hold285/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
Xhold296 hold296/I _7665_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
Xhold263 _7800_/Q hold263/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
Xhold274 hold274/I hold274/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
XFILLER_172_37 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_132_676 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_104_389 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_77_229 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_49_69 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_131_197 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_58_443 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7179_ _7393_/Q _7200_/A2 _7201_/B1 _7507_/Q _7200_/B1 _7387_/Q _7182_/A1 VDD VSS
+ gf180mcu_fd_sc_mcu7t5v0__aoi222_1
XFILLER_58_454 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_590 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_46_605 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2402 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_105_97 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_65_79 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_65_68 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_45_137 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1734 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1723 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1712 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_121_52 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1701 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_157_2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1767 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1756 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1745 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_81_490 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_54_693 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1778 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1789 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_167_551 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_81_89 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_10_741 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_139_286 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_108_673 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_122_153 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_77_785 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_37_605 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_92_744 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_64_435 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
Xinput9 mask_rev_in[14] input9/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_17_340 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3900_ _7813_/Q _6350_/A1 _6316_/A1 _7797_/Q _3901_/A4 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_4880_ _4448_/Z _4882_/A2 _4880_/B _7531_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_17_384 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_32_321 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3831_ hold123/Z _3787_/Z hold127/Z _3963_/A4 _3886_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand4_4
XFILLER_32_343 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6550_ hold504/Z _6553_/A2 _6551_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_3762_ _3762_/A1 _3762_/A2 _7974_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_20_527 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_20_549 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5501_ _5064_/B _5501_/A2 _5501_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__or2_1
XFILLER_72_2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3693_ _7378_/Q _3693_/ZN VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_145_201 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_145_212 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_145_223 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6481_ hold47/Z _6485_/A2 _6481_/B _7867_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_173_565 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_146_768 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_145_245 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5432_ _5778_/A1 _5162_/C _5686_/A2 _5725_/A1 _5435_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand4_1
X_5363_ _5600_/A1 _5363_/A2 _5797_/A1 _5363_/B _5703_/C VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai31_1
Xoutput335 _7949_/Q wb_dat_o[31] VDD VSS gf180mcu_fd_sc_mcu7t5v0__buf_8
Xoutput324 _7483_/Q wb_dat_o[21] VDD VSS gf180mcu_fd_sc_mcu7t5v0__buf_8
Xoutput302 _3927_/Z serial_data_2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__buf_8
Xoutput313 _7489_/Q wb_dat_o[11] VDD VSS gf180mcu_fd_sc_mcu7t5v0__buf_8
X_4314_ _4309_/S _4314_/A2 _4314_/B _7339_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_113_131 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7102_ _7827_/Q _7202_/A2 _7202_/B1 _7787_/Q _7763_/Q _7202_/C2 _7105_/A2 VDD VSS
+ gf180mcu_fd_sc_mcu7t5v0__aoi222_1
XFILLER_99_354 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5294_ _5212_/Z _5294_/A2 _5294_/B _5299_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_114_676 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_113_164 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_141_484 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_101_337 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7033_ _7695_/Q _7194_/A2 _7202_/B1 _7785_/Q _7035_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_68_741 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_19_28 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_4245_ _7724_/Q hold119/I _4594_/A1 _7401_/Q _4858_/A1 _7523_/Q _4248_/A2 VDD VSS
+ gf180mcu_fd_sc_mcu7t5v0__aoi222_2
XFILLER_28_605 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4176_ _7605_/Q _5920_/A1 _4219_/A2 input12/Z _4176_/C _4179_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi221_1
XFILLER_95_593 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_55_402 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_55_424 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7935_ _7935_/D _7961_/RN _7938_/CLK _7935_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XTAP_1019 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1008 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_7866_ _7866_/D _7901_/RN _7867_/CLK _7866_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_51_641 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_168_315 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6817_ _7682_/Q _6887_/B1 _6891_/B1 _7674_/Q _6819_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_23_354 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_51_674 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7797_ _7797_/D _7901_/RN _7797_/CLK _7797_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_11_538 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_149_562 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_137_702 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_6748_ _7639_/Q _6890_/A2 _6665_/Z _7743_/Q _6748_/C _6754_/B1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi221_1
XFILLER_176_392 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6679_ _7612_/Q _6647_/Z _6893_/B1 _7766_/Q _6681_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_151_215 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_151_248 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_2_247 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_160_771 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_120_602 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_78_516 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_120_646 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_104_197 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_59_763 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_86_582 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_86_571 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_73_210 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_59_785 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_18_104 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_19_638 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2210 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_100_392 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_74_744 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2243 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2232 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2221 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_132_95 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_92_33 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2287 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2276 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2265 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2254 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1542 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1531 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1520 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_14_321 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_2298 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1575 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1564 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1553 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_60 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_71 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_82 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_41_140 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1597 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1586 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_93 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_174_318 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_127_212 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_182_384 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_170_524 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_157_70 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_6_586 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_6_597 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_123_440 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_96_335 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_110_145 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_4030_ _4030_/A1 _4030_/A2 _4030_/A3 _4030_/A4 _4036_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand4_1
XFILLER_77_560 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_2_64 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_92_530 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5981_ hold41/Z _5987_/A2 _5981_/B hold319/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_4932_ _4906_/S _5210_/B _5138_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_7720_ _7720_/D _7901_/RN _7799_/CLK _7720_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_80_747 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_80_758 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_178_602 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7651_ _7651_/D _7961_/RN _7735_/CLK _7651_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_33_641 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_177_112 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_60_460 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4863_ _4863_/A1 _7285_/A2 _4867_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_32_173 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6602_ _6950_/A1 _6602_/A2 _7912_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_3814_ _3850_/A1 hold117/Z _3843_/A3 hold274/Z hold630/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand4_4
X_4794_ _7227_/I0 _7483_/Q _4795_/S _7483_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_32_184 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7582_ _7582_/D _7901_/RN _7582_/CLK _7582_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_158_392 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_158_370 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6533_ hold506/Z _6536_/A2 _6534_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_3745_ _4292_/B _4284_/A1 _7977_/Q _3747_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_21_18 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_173_351 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_119_768 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_6464_ hold47/Z _6468_/A2 _6464_/B _7859_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_173_362 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5415_ _5415_/A1 _5415_/A2 _5415_/B _5521_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_133_215 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3676_ _7606_/Q _7027_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_6395_ hold474/Z _6400_/A2 _6396_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_142_771 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xoutput176 _3698_/ZN mgmt_gpio_oeb[14] VDD VSS gf180mcu_fd_sc_mcu7t5v0__buf_8
X_5346_ _5692_/B _5692_/A2 _5347_/C VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_102_602 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xoutput198 _3678_/ZN mgmt_gpio_oeb[34] VDD VSS gf180mcu_fd_sc_mcu7t5v0__buf_8
Xoutput187 _3688_/ZN mgmt_gpio_oeb[24] VDD VSS gf180mcu_fd_sc_mcu7t5v0__buf_8
X_5277_ _5624_/A1 _5431_/B _5566_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_101_101 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_101_112 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_99_173 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7016_ _7016_/A1 _7016_/A2 _7016_/A3 _7016_/A4 _7026_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand4_1
XFILLER_87_357 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4228_ _7708_/Q _6141_/A1 _4759_/A1 _7468_/Q _4236_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_28_402 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_28_457 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_46_37 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4159_ _7621_/Q _5954_/A1 _4769_/A1 _7473_/Q _5971_/A1 _7629_/Q _4162_/A1 VDD VSS
+ gf180mcu_fd_sc_mcu7t5v0__aoi222_2
XFILLER_56_744 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_71_747 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_7918_ _7918_/D _7961_/RN _7940_/CLK _7918_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_43_438 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_43_449 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_102_76 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_7849_ _7849_/D _7901_/RN _7849_/CLK _7849_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_11_313 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_156_318 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_134_4 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_11_357 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_149_370 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_109_212 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_137_554 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_137_565 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_109_245 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_152_524 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_11_73 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_127_73 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_87_33 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_3_567 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_2_2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_132_292 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_94_806 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_120_498 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_143_83 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_47_744 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_47_799 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_2051 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2040 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_62_758 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_62_747 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_27_490 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_34_427 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_2095 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2084 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2073 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2062 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1350 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_15_641 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_159_134 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_1383 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1361 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1372 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_460 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1394 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
Xinput12 mask_rev_in[17] input12/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
Xinput45 mgmt_gpio_in[18] input45/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_168_91 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xinput34 mask_rev_in[8] input34/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
Xinput23 mask_rev_in[27] input23/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
Xinput56 mgmt_gpio_in[28] input56/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_116_738 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_115_215 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xinput89 spimemio_flash_io2_do input89/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
Xinput78 spi_csb input78/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
Xinput67 mgmt_gpio_in[3] input67/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_182_192 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_170_321 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_115_248 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5200_ _5230_/A1 _5663_/A1 _5200_/B _5202_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_6180_ _7726_/Q _6191_/A2 _6181_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_170_398 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5131_ _5006_/B _5344_/A2 _5480_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_35_2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5062_ _5006_/C _5616_/A1 _5062_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__and2_2
XFILLER_97_655 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_69_357 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_96_176 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4013_ _4013_/A1 _4013_/A2 _4013_/A3 _4013_/A4 _4013_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__and4_1
XFILLER_38_744 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_53_725 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_92_371 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_37_298 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_178_410 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_7703_ _7703_/D _7961_/RN _7735_/CLK _7703_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_80_566 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5964_ hold41/Z _5970_/A2 _5964_/B hold357/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_52_246 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4915_ _3728_/I _5369_/B _4915_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__and2_4
X_5895_ hold662/Z _5902_/A2 _5896_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_61_780 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_33_482 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_7634_ _7634_/D _7901_/RN _7820_/CLK _7634_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_166_605 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_139_808 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4846_ hold581/Z _4847_/A2 hold582/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_159_690 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_138_318 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7565_ _7565_/D input75/Z _7565_/CLK _7565_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
X_6516_ hold505/Z _6519_/A2 _6517_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_4777_ hold592/Z _4778_/A2 _4778_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_20_176 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_21_699 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3728_ _3728_/I _5338_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_8
XFILLER_174_660 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_106_204 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_7496_ _7496_/D _7912_/CLK _7496_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_3659_ _5195_/B _5011_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__inv_2
X_6447_ hold47/Z _6451_/A2 _6447_/B _7851_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_134_546 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_161_354 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6378_ hold421/Z _6383_/A2 _6379_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_115_771 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_88_600 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5329_ _5431_/B _5624_/A2 _5540_/C _5335_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_121_229 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_130_763 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_180_37 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_102_487 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_56_530 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_113_97 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_71_511 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_43_202 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_44_747 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_24_460 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_157_627 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_12_666 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_152_321 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_113_708 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_152_398 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_106_771 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_419 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_408 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_79_655 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_121_774 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_78_176 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_35_747 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_179_229 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_62_588 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_62_599 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_43_780 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_148_605 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5680_ _5680_/A1 _5779_/A2 _5680_/B1 _5680_/B2 _5680_/C _5681_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi221_1
X_4700_ _3819_/Z hold73/Z _4701_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_1
XTAP_1191 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1180 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_4631_ hold94/Z _3830_/Z _4631_/B hold95/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_30_463 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_147_159 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_128_351 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7350_ _7350_/D _7961_/RN _7353_/CLK _7350_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffsnq_2
X_4562_ hold578/Z _4563_/A2 _4563_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_7281_ _7520_/Q _7281_/A2 _7281_/B1 _7518_/Q _7519_/Q _7281_/C2 _7282_/A2 VDD VSS
+ gf180mcu_fd_sc_mcu7t5v0__aoi222_1
XFILLER_171_641 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_155_192 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xhold604 _7584_/Q hold604/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
X_6301_ _4448_/Z _6315_/A2 _6301_/B _7782_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_4493_ hold227/Z _4504_/A2 hold228/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
Xhold626 _7559_/Q hold626/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
Xhold615 _7374_/Q hold615/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
X_6232_ _4460_/Z _6242_/A2 _6232_/B hold125/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_143_354 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_131_505 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xhold659 _7521_/Q hold659/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
Xhold637 _7605_/Q hold637/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
Xhold648 _7397_/Q hold648/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
X_6163_ _7718_/Q _6174_/A2 _6164_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_920 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_931 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_942 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_953 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_5114_ _5648_/A1 _5058_/Z _5114_/A3 _5778_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand3_4
XFILLER_85_603 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6094_ _4454_/Z _6106_/A2 _6094_/B _7685_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
XTAP_964 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_975 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_986 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_5045_ _5538_/A1 _5042_/Z _5476_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_2
XFILLER_97_496 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_84_124 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_27_17 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_997 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_84_179 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_84_168 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_26_747 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_80_330 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6996_ _7669_/Q _7201_/B1 _7205_/A2 _7733_/Q _6997_/A4 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_5947_ hold41/Z _5953_/A2 _5947_/B hold457/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_41_739 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_80_396 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_179_785 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_178_273 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_139_638 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5878_ _4454_/Z _5880_/A2 _5878_/B _7584_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_7617_ _7617_/D _7901_/RN _7698_/CLK _7617_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
X_4829_ _7503_/Q _4828_/S _4830_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_119_373 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7548_ _7548_/D _7307_/Z _4418_/I1 _7548_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffnrnq_1
XFILLER_134_321 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7479_ _7479_/D _7944_/CLK _7479_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_161_184 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_134_398 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_88_430 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_68_46 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_130_571 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_103_785 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_88_463 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_76_625 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_356 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_48_316 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_124_52 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_84_34 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_75_146 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_29_552 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_90_116 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_90_105 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_44_544 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_140_73 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_25_780 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_32_739 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_44_599 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_252 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_241 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_230 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_157_424 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_285 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_274 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_263 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_129_115 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_12_463 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_296 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_172_416 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_145_619 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_8_456 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_153_641 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_144_129 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_180_460 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_152_151 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_180_471 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_165_70 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_3_150 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_79_430 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xhold1 hold1/I hold1/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
XFILLER_121_582 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_94_433 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_79_496 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_81_105 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_66_179 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6850_ _7433_/Q _7927_/Q _6850_/B _6852_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_62_330 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5801_ _5801_/A1 _5801_/A2 _5802_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_6781_ _7133_/S _6781_/A2 _6781_/B _7925_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_176_700 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3993_ _7689_/Q _6090_/A1 _5971_/A1 _7633_/Q _3993_/C _3999_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi221_4
X_5732_ _5732_/A1 _5732_/A2 _5732_/A3 _5732_/A4 _5795_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand4_1
XFILLER_176_744 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_175_232 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5663_ _5663_/A1 _5753_/A2 _5774_/B1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_31_783 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5594_ _4969_/C _5606_/B _5599_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_117_811 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7402_ _7402_/D _7961_/RN _7874_/CLK _7402_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
X_4614_ _4614_/A1 _7285_/A2 _4618_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_4545_ hold434/Z _4548_/A2 _4546_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_129_682 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_116_321 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xhold401 _7698_/Q hold401/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
X_7333_ input75/Z _4334_/Z _7333_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__and2_1
Xhold434 _7381_/Q hold434/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
XFILLER_144_663 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
Xhold412 _7681_/Q hold412/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
Xhold423 _7703_/Q hold423/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
Xhold445 _7679_/Q hold445/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
X_7264_ _7520_/Q _7264_/A2 _7266_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_171_460 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4476_ hold47/Z _4750_/I1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
Xhold467 _7844_/Q hold467/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
Xhold456 _7616_/Q hold456/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
Xhold478 hold478/I _7359_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
X_6215_ _4460_/Z _6225_/A2 _6215_/B hold243/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_131_357 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
Xhold489 _7351_/Q hold489/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
X_7195_ _7477_/Q _7195_/A2 _7195_/B1 _7471_/Q _7195_/C1 _7384_/Q _7198_/A2 VDD VSS
+ gf180mcu_fd_sc_mcu7t5v0__aoi222_1
X_6146_ _7710_/Q _6157_/A2 _6147_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_750 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_761 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_100_744 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_772 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_783 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_794 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_100_788 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_6077_ _4454_/Z _6089_/A2 _6077_/B _7677_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_46_809 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5028_ _5538_/A1 _5026_/Z _5545_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_85_499 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_72_116 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1916 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1905 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_54_37 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_1949 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1938 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1927 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_81_661 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_26_577 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_13_238 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_41_547 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6979_ _7002_/B _6979_/A2 _6979_/A3 _6979_/B _7931_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai31_1
XFILLER_179_593 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_70_58 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_154_405 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_135_630 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_5_415 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_135_641 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_107_354 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_102_2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_162_460 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_135_73 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_89_783 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_142 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_76_411 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_1_698 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_48_102 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_95_77 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_76_455 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_91_425 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_48_179 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_91_447 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_63_138 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_60_812 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_72_694 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_71_171 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_44_385 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_158_733 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_32_569 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_44_92 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_158_755 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_157_210 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_13_783 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_173_736 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_157_298 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_181_780 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_141_611 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_126_685 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_126_696 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_4330_ _4330_/I _7334_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_113_357 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_87_709 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4261_ _7347_/Q _4444_/A1 _5988_/A1 _7636_/Q _4262_/A4 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_140_176 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6000_ hold47/Z _6004_/A2 _6000_/B hold515/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_4192_ _7791_/Q _6316_/A1 _7285_/A1 _7961_/Q input21/Z _4239_/A2 _4194_/A3 VDD VSS
+ gf180mcu_fd_sc_mcu7t5v0__aoi222_1
XFILLER_95_753 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_39_135 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_7951_ _7951_/D _7959_/RN _4411_/I1 hold34/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_67_499 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_55_628 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_7882_ _7882_/D _7901_/RN _7890_/CLK _7882_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
X_6902_ _7912_/Q _7911_/Q _6936_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_4
X_6833_ _7853_/Q _6890_/B1 _6894_/C1 _7837_/Q _6834_/A4 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_50_300 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_51_812 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_50_333 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3976_ input40/Z _5903_/A1 _6209_/A1 _7745_/Q _3996_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_6764_ _7379_/Q _6882_/A2 _6894_/C1 _7834_/Q _6764_/C _6766_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi221_1
XFILLER_11_709 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_176_530 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5715_ _5408_/C _5715_/A2 _5715_/A3 _5732_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor3_1
X_6695_ _7733_/Q _6830_/B _6889_/A2 _7701_/Q _6767_/C _6697_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi221_1
X_5646_ _5510_/B _5646_/A2 _5646_/A3 _5740_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor3_1
XFILLER_136_405 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_164_747 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_108_118 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_163_246 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5577_ _5774_/A1 _4996_/Z _5062_/Z _5577_/B2 _5577_/C _5578_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi221_1
Xhold220 hold220/I _7667_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
XFILLER_117_641 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_151_419 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xhold242 _7742_/Q hold242/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
XFILLER_144_460 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xhold253 _7662_/Q hold253/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
XFILLER_116_151 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_2_418 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
Xhold231 _7365_/Q hold231/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
X_7316_ input75/Z _4334_/Z _7316_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__and2_1
X_4528_ hold709/Z _4531_/A2 _4529_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_7247_ _7247_/A1 _7280_/A2 _7277_/B _7247_/C _7248_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi211_1
X_4459_ hold5/Z _3810_/S hold6/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
Xhold286 _7796_/Q hold286/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
Xhold264 hold264/I _7800_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
Xhold275 hold630/I hold275/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
XFILLER_104_379 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
Xhold297 _7354_/Q hold297/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
XFILLER_131_187 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_131_176 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_86_742 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_58_411 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_7178_ _7178_/A1 _7178_/A2 _7178_/A3 _7184_/B1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor3_1
XFILLER_105_65 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6129_ hold209/Z _6140_/A2 hold210/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_580 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_591 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_73_425 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_73_414 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_58_499 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_45_105 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_1724 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1713 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1702 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_60_108 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_14_514 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_42_812 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1757 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1746 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1735 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_81_35 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_14_525 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1779 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1768 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_182_544 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_155_736 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_5_212 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_182_577 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_163_780 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_107_173 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_107_140 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_122_132 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_69_709 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_150_463 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_123_666 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_122_176 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_39_70 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_36_105 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_49_477 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_49_499 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xclkbuf_leaf_53_csclk clkbuf_3_6__f_csclk/Z _7694_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_36_127 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_36_149 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_33_801 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_33_812 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_45_672 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_51_119 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3830_ hold630/Z hold20/Z _3830_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__or2_4
Xclkbuf_leaf_68_csclk _7396_/CLK _7643_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_158_530 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3761_ _7974_/Q _3752_/I _3762_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_13_580 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_20_517 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5500_ _5064_/B _5501_/A2 _5641_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_146_758 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_146_747 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_118_449 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6480_ hold486/Z _6485_/A2 _6481_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_3692_ _7761_/Q _3692_/ZN VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_5431_ _5624_/A1 _5648_/B2 _5431_/B _5625_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_65_2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_161_739 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5362_ _5362_/A1 _5520_/C _5362_/B1 _5362_/B2 _7539_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_126_460 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xoutput325 _7484_/Q wb_dat_o[22] VDD VSS gf180mcu_fd_sc_mcu7t5v0__buf_8
Xoutput303 _4414_/Z serial_load VDD VSS gf180mcu_fd_sc_mcu7t5v0__buf_8
Xoutput314 _7490_/Q wb_dat_o[12] VDD VSS gf180mcu_fd_sc_mcu7t5v0__buf_8
X_4313_ _7339_/Q _4309_/S _4314_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_153_290 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7101_ _7819_/Q _7207_/A2 _7207_/B1 _7721_/Q _7101_/C _7105_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi221_1
XFILLER_113_121 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
Xoutput336 _7499_/Q wb_dat_o[3] VDD VSS gf180mcu_fd_sc_mcu7t5v0__buf_8
X_5293_ _5561_/B _5293_/A2 _5293_/A3 _5293_/A4 _5298_/A4 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand4_1
X_7032_ _7687_/Q _7189_/B1 _7188_/A2 _7378_/Q _7035_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_59_208 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_141_496 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_19_18 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4244_ _7612_/Q _5937_/A1 _4853_/A1 _7521_/Q _4244_/C _4248_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi221_2
XFILLER_67_241 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4175_ _7823_/Q _6384_/A1 _4614_/A1 _7410_/Q _4564_/A1 _7390_/Q _4179_/A1 VDD VSS
+ gf180mcu_fd_sc_mcu7t5v0__aoi222_1
XFILLER_83_712 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_82_200 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_27_105 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_55_436 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_83_778 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7934_ _7934_/D _7961_/RN _7938_/CLK _7934_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_24_801 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_36_672 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_42_108 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_1009 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_7865_ _7865_/D _7901_/RN _7865_/CLK _7865_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_51_631 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7796_ _7796_/D _7901_/RN _7799_/CLK _7796_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
X_6816_ _7626_/Q _6659_/Z _6884_/B1 _7690_/Q _6819_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_6747_ _6747_/A1 _6747_/A2 _6747_/A3 _6748_/C VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_50_174 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_149_574 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3959_ hold123/I _3787_/Z _3790_/Z _3963_/A4 _3959_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__or4_2
X_6678_ _7732_/Q _6830_/B _6893_/C1 _7628_/Q _6767_/C _6681_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi221_1
X_5629_ _5079_/Z _5433_/C _5629_/B _5684_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_145_780 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_4_6 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_132_463 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_78_506 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_2_259 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_116_75 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_104_176 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_116_86 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_93_509 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_2200 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_132_41 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_46_458 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2244 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2233 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2222 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2211 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_73_266 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_15_812 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2277 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2266 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2255 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1532 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1521 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1510 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_61_428 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_27_683 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_54_491 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2299 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2288 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1576 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1565 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1554 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1543 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_50 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_61 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_72 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_83 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_1598 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1587 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_94 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_128_747 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_128_736 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_182_352 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_182_341 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_128_769 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_127_246 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_41_93 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_143_739 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_108_460 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_51_8 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_135_290 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_173_70 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_151_783 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_150_282 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_123_496 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_111_636 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_110_102 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_69_539 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_110_179 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_65_712 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_37_425 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5980_ hold318/Z _5987_/A2 _5981_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_92_553 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_64_266 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_24_108 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_4931_ _5302_/A1 _5195_/B _5210_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__or2_1
XFILLER_80_737 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_17_160 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4862_ _4454_/Z _4862_/A2 _4862_/B _7524_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_7650_ _7650_/D _7961_/RN _7650_/CLK _7650_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
X_3813_ _3810_/S hold273/Z hold274/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_4
XFILLER_20_314 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6601_ _7912_/Q _6618_/A3 _6601_/B _6602_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_177_179 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_165_319 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4793_ _4807_/A1 _4795_/S _4793_/B _7482_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_7581_ _7581_/D _7961_/RN _7961_/CLK _7581_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_118_202 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6532_ hold47/Z _6536_/A2 _6532_/B _7891_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_3744_ _3744_/A1 _3751_/A2 _4284_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_4
XFILLER_173_341 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6463_ hold516/Z _6468_/A2 _6464_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_3675_ _7605_/Q _6707_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_161_503 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_134_739 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_134_717 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_127_780 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5414_ _5414_/A1 _5414_/A2 _5414_/A3 _5414_/A4 _5415_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor4_1
X_6394_ hold41/Z _6400_/A2 _6394_/B _7826_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
Xoutput177 _3697_/ZN mgmt_gpio_oeb[15] VDD VSS gf180mcu_fd_sc_mcu7t5v0__buf_8
X_5345_ _5176_/B _5573_/A1 _5477_/B2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_114_463 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_99_152 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_99_141 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_88_804 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xoutput199 _4393_/ZN mgmt_gpio_oeb[35] VDD VSS gf180mcu_fd_sc_mcu7t5v0__buf_8
Xoutput188 _3687_/ZN mgmt_gpio_oeb[25] VDD VSS gf180mcu_fd_sc_mcu7t5v0__buf_8
XFILLER_102_636 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5276_ _5409_/B2 _5350_/A3 _5412_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_87_336 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7015_ _7872_/Q _7195_/C1 _7015_/B _7016_/A4 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_4227_ _7668_/Q _6056_/A1 _5846_/A1 _7571_/Q _4240_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_55_233 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4158_ _4158_/A1 _4158_/A2 _4158_/A3 _4158_/A4 _4204_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand4_2
XFILLER_56_756 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4089_ input54/Z _5886_/A1 _5971_/A1 _7630_/Q _4090_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_16_609 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_28_469 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_102_33 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_70_225 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_43_428 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7917_ _7917_/D _7961_/RN _7940_/CLK _7917_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_70_247 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_62_37 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_24_664 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_178_37 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_168_135 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_168_124 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7848_ _7848_/D _7901_/RN _7849_/CLK _7848_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffsnq_1
XFILLER_23_152 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_23_141 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7779_ _7779_/D _7901_/RN _7851_/CLK _7779_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_51_494 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_168_179 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_109_202 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_137_544 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_125_706 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_180_812 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_125_728 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_152_558 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_133_783 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_105_496 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_47_712 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_143_73 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_74_531 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_19_425 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_19_469 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_2052 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2041 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2030 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2085 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2074 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2063 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1340 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_15_631 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_2096 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1384 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1362 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1373 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1351 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_15_697 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_42_450 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_159_168 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_1395 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_174_105 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xinput13 mask_rev_in[18] input13/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
Xinput46 mgmt_gpio_in[19] input46/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_174_138 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_168_81 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_168_70 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
Xinput35 mask_rev_in[9] input35/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
Xinput24 mask_rev_in[28] input24/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_171_812 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_155_363 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
Xinput57 mgmt_gpio_in[29] input57/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
Xinput79 spi_enabled _4396_/S VDD VSS gf180mcu_fd_sc_mcu7t5v0__buf_2
Xinput68 mgmt_gpio_in[5] input68/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_115_238 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_109_780 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_131_709 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_124_761 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5130_ _5735_/A2 _5179_/B _5749_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_69_325 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5061_ _3722_/I _3723_/I _5006_/B _5616_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor3_4
XFILLER_28_2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4012_ _7712_/Q _6141_/A1 hold119/I _7728_/Q _4013_/A4 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_111_499 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_80_501 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_53_704 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xclkbuf_3_6__f_csclk clkbuf_0_csclk/Z clkbuf_3_6__f_csclk/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_80_534 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_80_523 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_65_586 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5963_ hold356/Z _5970_/A2 _5964_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_25_428 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_37_277 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4914_ _4914_/A1 _4914_/A2 _4914_/A3 _4914_/A4 _4914_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__or4_2
X_7702_ _7702_/D _7961_/RN _7702_/CLK _7702_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffsnq_1
XFILLER_52_236 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5894_ hold73/Z _5902_/A2 _5894_/B _7591_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_7633_ _7633_/D _7901_/RN _7812_/CLK _7633_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_60_280 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4845_ _4448_/Z _4847_/A2 _4845_/B _7507_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_21_645 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_32_29 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_33_494 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_148_29 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_7564_ _7564_/D input75/Z _7565_/CLK _7564_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffsnq_2
X_4776_ _4448_/Z _4778_/A2 _4776_/B _7474_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_3727_ _3727_/I _5201_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__inv_8
X_6515_ hold47/Z _6519_/A2 _6515_/B _7883_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_180_108 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_174_672 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_162_812 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7495_ _7495_/D _7961_/RN _7627_/CLK _7495_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
X_3658_ _3658_/I _7282_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_6446_ hold472/Z _6451_/A2 _6447_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_6377_ hold41/Z _6383_/A2 _6377_/B _7818_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_121_208 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5328_ _5333_/A3 _5495_/B2 _5540_/C VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_2
XFILLER_115_783 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_527 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_87_144 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_76_807 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5259_ _4996_/Z _5087_/B _5433_/C _5701_/C VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand3_2
XFILLER_29_712 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_57_59 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_28_266 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_44_715 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_71_567 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_51_280 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_169_499 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_169_488 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_156_105 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_132_2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_12_656 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_11_144 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_8_605 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_156_149 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_153_812 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_164_171 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_138_84 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_3_310 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_3_354 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_3_376 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_409 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_154_61 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_154_83 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_120_274 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_93_136 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_35_704 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_47_81 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_170_93 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_90_810 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_62_534 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_47_586 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_34_236 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_34_247 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_62_578 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1192 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1181 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1170 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_179_91 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_175_425 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4630_ _3830_/Z _4460_/Z _4631_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_162_119 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_162_108 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_144_812 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6300_ hold740/Z _6315_/A2 _6301_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_4561_ _4448_/Z _4563_/A2 _4561_/B _7387_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_7280_ _4376_/B _7280_/A2 _7280_/A3 _7282_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand3_1
Xhold627 _7463_/Q hold627/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
XFILLER_143_300 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
Xhold605 _7799_/Q hold605/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
XFILLER_116_547 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_7_682 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_4492_ _4454_/Z _4504_/A2 _4492_/B hold700/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
Xhold616 _7394_/Q hold616/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
X_6231_ _7750_/Q _6242_/A2 _6232_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
Xhold638 _7708_/Q hold638/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
Xhold649 _7621_/Q hold649/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
XFILLER_143_388 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6162_ _4454_/Z _6174_/A2 _6162_/B _7717_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
XTAP_910 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_5113_ _5496_/A1 _5458_/C _5661_/A1 _5473_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor3_1
XFILLER_112_731 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_69_144 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_921 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_932 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_943 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_6093_ hold713/Z _6106_/A2 _6094_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_954 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_965 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_976 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_987 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_5044_ _5452_/C _5543_/C _5475_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_111_296 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_998 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_38_575 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_53_567 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6995_ _7815_/Q _7207_/A2 _7207_/B1 _7717_/Q _7205_/B1 _7741_/Q _6997_/A3 VDD VSS
+ gf180mcu_fd_sc_mcu7t5v0__aoi222_1
X_5946_ hold456/Z _5953_/A2 _5947_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_53_578 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_159_39 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5877_ hold604/Z _5880_/A2 _5878_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_43_39 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_166_425 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_166_403 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_138_105 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7616_ _7616_/D _7961_/RN _7704_/CLK _7616_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
X_4828_ _7228_/I0 _7502_/Q _4828_/S _7502_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_181_428 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_135_812 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_119_363 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_5_619 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4759_ _4759_/A1 _7285_/A2 _4763_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_7547_ _7547_/D _7901_/RN _7582_/CLK _7547_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_4_129 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_7478_ _7478_/D _7944_/CLK _7478_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_162_653 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_161_130 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_161_141 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6429_ hold519/Z _6434_/A2 _6430_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_104_6 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_76_615 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_76_637 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_48_328 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_84_46 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_84_24 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_75_169 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_16_203 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_16_247 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_17_73 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_44_534 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_242 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_231 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_220 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_71_386 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_31_239 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_169_274 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_286 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_275 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_264 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_253 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_297 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_144_108 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_138_661 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_138_672 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_126_812 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_152_130 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_141_804 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_165_82 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_140_314 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xhold2 hold2/I hold2/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
XFILLER_66_125 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_181_70 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_35_534 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3992_ _3992_/A1 _3992_/A2 _3992_/A3 _3993_/C VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand3_1
X_5800_ _5800_/A1 _5800_/A2 _5801_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_90_673 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6780_ _7925_/Q _7133_/S _6781_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_22_206 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_35_567 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5731_ _5104_/B _5608_/B _5731_/B _5732_/A4 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_95_2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_176_767 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5662_ _5662_/A1 _5797_/A2 _5774_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_30_250 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_31_773 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5593_ _5608_/A1 _5167_/B _5606_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__or2_2
X_4613_ _4454_/Z _4613_/A2 _4613_/B _7408_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_7401_ _7401_/D _7961_/RN _7756_/CLK _7401_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
X_4544_ hold47/Z _4548_/A2 _4544_/B _7380_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_163_428 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
Xhold402 _7618_/Q hold402/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
X_7332_ input75/Z _4334_/Z _7332_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__and2_1
X_7263_ _7263_/A1 _7277_/B _7263_/B _7954_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_143_141 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xhold435 _7666_/Q hold435/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
XFILLER_128_193 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
Xhold424 _7671_/Q hold424/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
Xhold413 _7609_/Q hold413/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
X_4475_ _7970_/Q _7506_/Q hold46/Z hold47/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_4
X_6214_ hold242/Z _6225_/A2 _6215_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
Xhold446 _7736_/Q hold446/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
Xhold468 _7763_/Q hold468/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
XFILLER_89_206 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xhold457 hold457/I _7616_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
XFILLER_143_185 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
Xhold479 _7779_/Q hold479/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
XFILLER_98_740 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_7194_ _7524_/Q _7194_/A2 _7194_/B1 _7505_/Q _7194_/C1 _7410_/Q _7199_/A2 VDD VSS
+ gf180mcu_fd_sc_mcu7t5v0__aoi222_1
X_6145_ _4454_/Z _6157_/A2 _6145_/B _7709_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
XTAP_740 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_751 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_100_734 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_97_294 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_97_272 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_97_283 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6076_ hold689/Z _6089_/A2 _6077_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_762 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_773 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_784 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_795 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_5027_ _5538_/A1 _5026_/Z _5027_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__and2_1
XTAP_1906 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_81_651 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_26_534 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1939 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1928 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1917 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_110_33 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_13_228 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6978_ _7604_/Q _6949_/I _6979_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_167_712 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_110_77 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5929_ hold441/Z _5936_/A2 _5930_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_166_211 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_139_425 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_70_37 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_21_272 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_126_108 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_108_812 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_21_283 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_182_737 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_181_247 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_134_130 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_150_601 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_134_152 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_79_57 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_122_347 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_122_336 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_88_250 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_135_85 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_76_445 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_91_415 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_76_489 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_29_372 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_29_361 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_151_73 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_17_567 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_9_700 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_12_250 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_9_722 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_145_428 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_67_6 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_60_92 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_8_276 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_172_247 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_160_409 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_125_141 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_125_196 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_113_347 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_5_98 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4260_ _4260_/A1 _4260_/A2 _4260_/A3 _4260_/A4 _4263_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand4_1
XFILLER_101_509 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_4191_ _7396_/Q _4579_/A1 _4774_/A1 _7475_/Q _4194_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_79_294 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_79_283 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_67_423 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_10_2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_7950_ _7950_/D _7959_/RN _4411_/I1 hold14/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_82_415 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_36_810 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7881_ _7881_/D _7901_/RN _7881_/CLK _7881_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
X_6901_ _7931_/Q _7133_/S _6979_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_6832_ _7845_/Q _6894_/A2 _6659_/Z _7627_/Q _6834_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_90_492 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_149_712 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3975_ _7771_/Q _6265_/A1 _6418_/A1 _7843_/Q _3996_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_6763_ _6763_/A1 _6763_/A2 _6763_/A3 _6764_/C VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_50_345 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_148_211 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5714_ _5714_/A1 _5099_/B _5714_/B1 _5722_/A1 _5715_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai22_1
XFILLER_31_570 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_50_389 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6694_ _7839_/Q _6894_/A2 _6659_/Z _7621_/Q _6697_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_5645_ _5645_/A1 _5687_/B _5645_/A3 _5099_/B _5741_/A3 _5646_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai32_1
XFILLER_108_108 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5576_ _4960_/Z _5663_/A1 _5372_/Z _5576_/B2 _5576_/C _5715_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai221_1
XFILLER_156_29 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_129_491 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xhold210 hold210/I _6130_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
Xhold243 hold243/I _7742_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
Xhold221 _7635_/Q hold221/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
X_7315_ _7901_/RN _4334_/Z _7315_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__and2_1
Xhold232 hold232/I _4511_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
X_4527_ _4527_/A1 _7285_/A2 _4531_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_7246_ _7246_/A1 _7246_/A2 _7247_/C VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_4458_ _7506_/Q hold28/Z hold29/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
Xhold287 hold287/I _6330_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
Xhold254 hold254/I _7662_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
Xhold276 hold276/I hold276/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
XFILLER_131_122 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
Xhold265 _7824_/Q hold265/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
XFILLER_132_678 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_131_144 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_32
Xhold298 hold298/I _4487_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
XFILLER_49_49 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_7177_ _7177_/A1 _7177_/A2 _7177_/A3 _7177_/A4 _7178_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand4_1
XFILLER_105_33 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4389_ _4387_/S _7897_/Q _4389_/B _4389_/ZN VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_2
X_6128_ _4454_/Z _6140_/A2 _6128_/B _7701_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
XTAP_570 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_100_531 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_58_467 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_581 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_592 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_85_286 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6059_ hold725/Z _6072_/A2 _6060_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_26_331 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1725 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1714 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1703 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1758 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1747 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1736 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_121_54 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_81_25 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_26_386 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_54_695 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1769 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_139_200 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_14_41 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_22_581 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_182_534 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_182_523 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_127_428 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_6_725 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_154_247 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_6_747 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_142_409 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_30_51 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_146_73 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_122_100 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_1_441 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_89_570 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_103_380 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_1_496 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_49_467 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_162_94 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_18_810 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_36_117 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_91_212 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_64_459 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_17_353 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_32_312 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_177_317 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3760_ _3760_/A1 _3756_/B _3765_/A2 _3760_/B2 _7975_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_60_676 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_13_570 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_32_389 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5430_ _5247_/B _5724_/B _5550_/B _5725_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_3691_ _7769_/Q _3691_/ZN VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_173_567 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_161_729 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_5361_ _5361_/A1 _5361_/A2 _5362_/B2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_126_450 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
Xoutput326 _7485_/Q wb_dat_o[23] VDD VSS gf180mcu_fd_sc_mcu7t5v0__buf_8
Xoutput304 _4413_/Z serial_resetn VDD VSS gf180mcu_fd_sc_mcu7t5v0__buf_8
Xoutput315 _7491_/Q wb_dat_o[13] VDD VSS gf180mcu_fd_sc_mcu7t5v0__buf_8
XFILLER_58_2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4312_ _7338_/Q _7414_/Q _4312_/B _4314_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_7100_ _7100_/A1 _7100_/A2 _7100_/A3 _7101_/C VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand3_1
X_5292_ _5724_/B _5624_/B _5292_/B _5293_/A4 VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_5_780 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xoutput337 _7500_/Q wb_dat_o[4] VDD VSS gf180mcu_fd_sc_mcu7t5v0__buf_8
XFILLER_114_678 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_113_144 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_102_807 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_7031_ _7801_/Q _7191_/B1 _7194_/C1 _7809_/Q _7035_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_4243_ _4243_/A1 _4243_/A2 _4243_/A3 _4244_/C VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_68_765 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_67_231 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_4174_ _4174_/A1 _4174_/A2 _4174_/A3 _4174_/A4 _4187_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand4_1
XFILLER_67_286 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7933_ _7933_/D _7961_/RN _7938_/CLK _7933_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_82_267 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_36_640 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7864_ _7864_/D _7901_/RN _7867_/CLK _7864_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffsnq_1
XFILLER_63_492 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6815_ _6815_/A1 _6815_/A2 _6815_/A3 _6815_/A4 _6825_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand4_1
X_7795_ _7795_/D _7901_/RN _7799_/CLK _7795_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
X_6746_ _7849_/Q _6890_/B1 _6894_/C1 _7833_/Q _6747_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_3958_ _3958_/A1 _4427_/B _3958_/B1 _3958_/B2 _7554_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_164_523 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_109_428 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3889_ _7627_/Q _5954_/A1 _4505_/A1 _7370_/Q _3892_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_6677_ _6677_/A1 _6677_/A2 _6677_/A3 _6677_/A4 _6684_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand4_1
XFILLER_164_534 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_5628_ _5363_/B _5627_/Z _5634_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_5559_ _5559_/A1 _5415_/B _5560_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_3_706 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_132_453 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_104_188 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7229_ _7949_/Q _7228_/S _7230_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_2201 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_74_757 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_73_212 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2234 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2223 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2212 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2278 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2267 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2256 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2245 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_162_2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1533 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1522 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1511 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1500 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_92_46 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_40 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_2289 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1566 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1555 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1544 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_14_345 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_51 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_62 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_73 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_42_632 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1599 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1588 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1577 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_25_73 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_84 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_42_676 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_95 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_167_361 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_155_523 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_182_331 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_155_567 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_10_584 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_10_573 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_157_94 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_6_588 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_69_507 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_150_272 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_150_250 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_96_315 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_2_44 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_49_231 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_49_286 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_52_407 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_4930_ _5195_/B _5201_/B _5210_/A3 _4926_/Z _4930_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__or4_4
XFILLER_18_673 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4861_ hold672/Z _4862_/A2 _4862_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_178_637 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3812_ hold272/Z _3799_/B _7414_/Q _3812_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_33_676 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6600_ _7434_/Q _6599_/Z _6601_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_4792_ _7482_/Q _4795_/S _4793_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_7580_ _7580_/D _7961_/RN _7580_/CLK _7580_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_2
XFILLER_20_337 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_6531_ hold522/Z _6536_/A2 _6532_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_3743_ _7346_/Q _7345_/Q _7344_/Q _4206_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor3_4
X_3674_ hold88/Z _7278_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_146_534 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_118_247 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6462_ hold41/Z _6468_/A2 _6462_/B _7858_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_146_578 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_118_269 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5413_ _5732_/A1 _5413_/A2 _5413_/A3 _5588_/A3 _5414_/A4 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand4_1
X_6393_ hold411/Z _6400_/A2 _6394_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_5344_ _5344_/A1 _5344_/A2 _5623_/A1 _5350_/A3 _5545_/A2 _5687_/B _5347_/B VDD VSS
+ gf180mcu_fd_sc_mcu7t5v0__oai33_1
XFILLER_114_453 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_709 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
Xoutput167 _4431_/Z debug_in VDD VSS gf180mcu_fd_sc_mcu7t5v0__buf_8
Xoutput178 _3696_/ZN mgmt_gpio_oeb[16] VDD VSS gf180mcu_fd_sc_mcu7t5v0__buf_8
Xoutput189 _3686_/ZN mgmt_gpio_oeb[26] VDD VSS gf180mcu_fd_sc_mcu7t5v0__buf_8
X_5275_ _5714_/B1 _5623_/A1 _5712_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_141_283 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7014_ _7014_/A1 _7014_/A2 _7015_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_4226_ _7558_/Q _5817_/A1 _4522_/A1 _7371_/Q _4267_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_101_169 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4157_ _7661_/Q _6039_/A1 _6333_/A1 _7799_/Q _4158_/A4 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_56_713 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_55_212 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_83_565 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4088_ _7349_/Q _4444_/A1 _4249_/A2 input26/Z _4505_/A1 _7365_/Q _4090_/A2 VDD VSS
+ gf180mcu_fd_sc_mcu7t5v0__aoi222_2
X_7916_ _7916_/D _7961_/RN _7938_/CLK _7916_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
X_7847_ _7847_/D _7901_/RN _7851_/CLK _7847_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffsnq_1
XFILLER_169_637 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_24_676 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_51_451 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_7778_ _7778_/D _7901_/RN _7853_/CLK _7778_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
X_6729_ _6729_/A1 _6729_/A2 _6729_/A3 _6728_/Z _6731_/B1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand4_1
XFILLER_164_331 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_109_225 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_137_567 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xclkbuf_leaf_52_csclk clkbuf_3_6__f_csclk/Z _7735_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_87_13 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_3_558 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_132_250 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_87_68 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
Xclkbuf_leaf_67_csclk _7396_/CLK _7645_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_143_63 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_59_551 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_86_392 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_59_595 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_2042 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2020 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2031 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_74_598 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_61_215 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_2086 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2075 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2064 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2053 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1341 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1330 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2097 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1363 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1374 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1352 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_30_602 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1396 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1385 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_128_534 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xinput14 mask_rev_in[19] input14/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
Xinput25 mask_rev_in[29] input25/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
Xinput36 mgmt_gpio_in[0] input36/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
Xinput69 mgmt_gpio_in[6] input69/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_10_392 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
Xinput47 mgmt_gpio_in[1] input47/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
Xinput58 mgmt_gpio_in[2] input58/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__buf_3
XFILLER_109_792 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_97_602 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_170_389 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_151_570 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_123_272 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5060_ _5319_/C _5692_/B _5301_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_123_283 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_96_134 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_69_348 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_84_318 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4011_ _7736_/Q _6192_/A1 _6090_/A1 _7688_/Q _4013_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_37_212 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5962_ hold73/Z _5970_/A2 _5962_/B hold528/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_4913_ _4914_/A1 _4914_/A2 _4914_/A3 _4914_/A4 _5211_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor4_4
X_7701_ _7701_/D _7961_/RN _7701_/CLK _7701_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffsnq_1
X_5893_ hold363/Z _5902_/A2 _5894_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_7632_ _7632_/D _7901_/RN _7820_/CLK _7632_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_60_270 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4844_ hold666/Z _4847_/A2 _4845_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_4775_ hold677/Z _4778_/A2 _4776_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_7563_ _7563_/D input75/Z _7567_/CLK _7563_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
X_3726_ _5199_/B _5200_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__inv_8
XFILLER_119_534 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6514_ hold524/Z _6519_/A2 _6515_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_146_342 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_119_567 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_107_707 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7494_ _7494_/D _7961_/RN _7532_/CLK _7494_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
X_6445_ hold41/Z _6451_/A2 _6445_/B _7850_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_3657_ _7916_/Q _6905_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_2
X_6376_ hold444/Z _6383_/A2 _6377_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_114_250 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5327_ _5431_/B _5624_/A2 _5803_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_88_602 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5258_ _5290_/B _5409_/B2 _5258_/B _5585_/C VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_5189_ _5658_/B _5643_/A2 _5642_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_68_392 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4209_ _4075_/B hold107/Z _5846_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_28_212 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_29_779 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_43_215 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_71_557 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_71_546 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_71_535 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_169_434 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_12_602 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_12_646 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_11_101 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_24_473 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_169_478 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_125_2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_180_621 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_164_183 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_98_34 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_180_676 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_152_334 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_152_389 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_133_570 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_112_209 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_79_624 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_3_366 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_105_283 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_67_808 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_94_605 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_66_318 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_66_307 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_19_212 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_170_50 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_47_543 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_47_565 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_28_790 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_50_708 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_63_70 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_179_70 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1182 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1171 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1160 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_63_92 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_30_410 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_42_270 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1193 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_147_139 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_8_65 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4560_ hold678/Z _4563_/A2 _4561_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_156_662 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_156_684 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_116_526 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_116_515 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
Xhold606 _7532_/Q hold606/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
X_4491_ hold698/Z _4504_/A2 hold699/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
Xhold617 _7467_/Q hold617/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
X_6230_ _4454_/Z _6242_/A2 _6230_/B _7749_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
Xhold628 _7340_/Q hold628/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
Xhold639 _7863_/Q hold639/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
X_6161_ hold608/Z _6174_/A2 _6162_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_40_2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_900 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_112_743 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5112_ _4996_/Z _5793_/A2 _5673_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_97_432 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_911 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_922 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_933 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_944 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_111_242 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6092_ _4448_/Z _6106_/A2 _6092_/B _7684_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
XTAP_955 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_966 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_977 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_5043_ _5548_/A1 _5043_/A2 _5543_/C VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_4
XFILLER_111_286 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_85_638 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_988 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_999 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
Xclkbuf_0_wbbd_sck _7958_/Q clkbuf_0_wbbd_sck/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_93_671 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_25_215 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_26_738 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_92_192 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_80_321 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6994_ _7879_/Q _7203_/B1 _7204_/A2 _7839_/Q _6997_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_5945_ hold73/Z _5953_/A2 _5945_/B hold547/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_80_376 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_43_29 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5876_ _4460_/Z _5880_/A2 _5876_/B hold33/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_33_281 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_139_618 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_7615_ _7615_/D _7961_/RN _7704_/CLK _7615_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffsnq_1
X_4827_ _7227_/I0 _7501_/Q _4828_/S _7501_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_21_465 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_135_802 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4758_ _4454_/Z _4758_/A2 _4758_/B _7467_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_7546_ _7546_/D _7901_/RN _7582_/CLK _7546_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
X_4689_ hold164/Z _3819_/Z _4689_/B hold165/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_4_108 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7477_ _7477_/D _7961_/RN _7572_/CLK _7477_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
X_3709_ _7631_/Q _3709_/ZN VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_108_33 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6428_ hold41/Z _6434_/A2 _6428_/B _7842_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_162_676 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_134_389 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_115_570 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6359_ hold320/Z _6366_/A2 _6360_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_103_732 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_68_37 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_314 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_102_242 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_76_605 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_75_126 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_29_510 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_48_318 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_56_362 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_17_749 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XPHY_210 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_25_771 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_243 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_232 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_221 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_24_270 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_31_229 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_276 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_265 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_254 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_12_443 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_169_286 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_298 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_287 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_33_73 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_40_796 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_149_95 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_149_73 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_153_621 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_152_120 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_99_708 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_113_518 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_113_529 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_113_507 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_3_141 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_180_495 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
Xhold3 hold3/I hold3/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
XFILLER_67_638 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_66_104 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_94_479 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_47_373 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_62_321 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3991_ _7665_/Q _6039_/A1 _6192_/A1 _7737_/Q _3992_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_50_505 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5730_ _5763_/A3 _5730_/A2 _5738_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_16_782 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_50_538 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_50_527 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_175_212 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5661_ _5661_/A1 _5661_/A2 _5661_/B _5774_/C VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_88_2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_31_796 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_7400_ _7400_/D _7961_/RN _7756_/CLK _7400_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_135_109 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_5592_ _5608_/A1 _5167_/B _5753_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_4612_ hold576/Z _4613_/A2 _4613_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_4543_ hold473/Z _4548_/A2 _4544_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_7331_ input75/Z _4334_/Z _7331_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__and2_1
X_7262_ _7262_/A1 _7280_/A2 _7277_/B _7262_/C _7263_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi211_1
Xhold436 hold436/I _7666_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
Xhold414 _7737_/Q hold414/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
Xhold425 hold425/I _7671_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
Xhold403 hold403/I _7618_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
X_4474_ _7506_/Q _7268_/A1 hold46/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_144_676 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
Xhold458 _7868_/Q hold458/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
XFILLER_116_389 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xhold469 _7869_/Q hold469/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
Xhold447 _7789_/Q hold447/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
X_6213_ _4454_/Z _6225_/A2 _6213_/B _7741_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_7193_ _7396_/Q _7193_/A2 _7193_/B1 _7473_/Q _7193_/C1 _7532_/Q _7199_/A1 VDD VSS
+ gf180mcu_fd_sc_mcu7t5v0__aoi222_1
X_6144_ hold565/Z _6157_/A2 _6145_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_131_359 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_58_616 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_58_605 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_730 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_741 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_752 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_6075_ _4448_/Z _6089_/A2 _6075_/B _7676_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_100_724 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_98_796 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_763 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_774 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_38_29 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_785 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_5026_ _5548_/A1 _5535_/A1 _5026_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__and2_1
XTAP_796 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_66_682 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_54_811 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1907 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_81_641 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1929 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1918 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_6977_ _7210_/A2 _6977_/A2 _6977_/A3 _6977_/A4 _6979_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor4_1
XFILLER_14_719 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_53_354 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5928_ hold73/Z _5936_/A2 _5928_/B _7607_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_110_67 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_22_741 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5859_ hold381/Z _5868_/A2 _5860_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_182_727 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_181_226 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_181_215 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_107_312 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_5_428 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7529_ _7529_/D _7961_/RN _7960_/CLK _7529_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_135_632 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_134_120 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_79_36 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_107_367 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_150_657 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_135_20 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_111 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_89_774 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_89_763 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_89_785 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_177 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_49_638 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_130_392 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_95_68 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_88_295 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_76_479 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_44_321 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_151_96 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_17_557 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_157_212 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_81_9 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_9_712 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_176_60 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_125_120 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_126_676 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_99_527 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_153_495 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_113_337 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_5_88 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4190_ _7783_/Q _6299_/A1 _6418_/A1 _7839_/Q _7580_/Q hold26/I _4194_/A1 VDD VSS
+ gf180mcu_fd_sc_mcu7t5v0__aoi222_1
XFILLER_67_446 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_39_126 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_7880_ _7880_/D _7901_/RN _7893_/CLK _7880_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffsnq_1
XFILLER_63_641 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_63_630 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6900_ _7133_/S _6900_/A2 _6900_/B _7930_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_6831_ _7707_/Q _6889_/A2 _6834_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_35_354 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_90_471 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_35_376 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3974_ _7657_/Q _6022_/A1 hold134/I _7819_/Q _3989_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_6762_ _7664_/Q _6885_/A2 _6893_/B1 _7770_/Q _6763_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_62_195 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_176_510 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5713_ _5716_/A1 _5716_/A2 _5716_/A3 _5795_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand3_1
X_6693_ _7613_/Q _6647_/Z _6887_/B1 _7677_/Q _6705_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_50_368 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_50_379 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_136_407 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5644_ _5644_/A1 _5644_/A2 _5644_/A3 _5804_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_164_738 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_163_204 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_163_215 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5575_ _5212_/Z _5575_/A2 _5768_/A3 _5576_/C VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_163_248 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_116_120 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xhold200 _7654_/Q hold200/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
Xhold211 hold211/I _7702_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
X_7314_ input75/Z _4334_/Z _7314_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__and2_1
Xhold244 _7848_/Q hold244/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
Xhold222 hold222/I _7635_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
Xhold233 hold233/I _7365_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
X_4526_ _4454_/Z _4526_/A2 _4526_/B _7372_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_7245_ _7520_/Q _7245_/A2 _7245_/B1 _7519_/Q _7246_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_171_292 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xhold255 _7464_/Q hold255/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
Xhold277 _7722_/Q hold277/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
XFILLER_132_646 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
Xhold266 hold266/I _6390_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
XFILLER_104_337 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4457_ hold246/Z _4487_/A1 hold247/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
Xhold288 hold288/I _7796_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
Xhold299 hold299/I _7354_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
X_7176_ _7391_/Q _6938_/I _7188_/A2 _7756_/Q _7177_/A4 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_4388_ _4387_/S input92/Z _4389_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_6127_ hold721/Z _6140_/A2 _6128_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_560 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_112_392 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_86_744 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_571 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_582 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_593 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_85_276 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_6058_ _4448_/Z _6072_/A2 _6058_/B _7668_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_5009_ _5199_/B _4898_/Z _4915_/Z _5005_/Z _5529_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand4_4
XFILLER_26_321 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_164_6 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1715 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_121_44 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_1704 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_26_343 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1748 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1737 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1726 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_14_538 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_14_516 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1759 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_41_357 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_179_370 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_139_212 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_167_565 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_10_733 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_155_727 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_30_41 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_108_676 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_107_164 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_123_668 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_122_145 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_110_318 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_162_84 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_77_777 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_92_747 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_91_235 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_91_246 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_45_641 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_45_674 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_60_666 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_158_598 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_158_587 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_158_576 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_146_749 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_145_215 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_3690_ _7777_/Q _3690_/ZN VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_161_708 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_145_237 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_5360_ _5415_/B _5360_/A2 _5360_/B _7279_/B _5361_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_114_602 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xoutput305 _4430_/Z spi_sdi VDD VSS gf180mcu_fd_sc_mcu7t5v0__buf_8
Xoutput316 _7492_/Q wb_dat_o[14] VDD VSS gf180mcu_fd_sc_mcu7t5v0__buf_8
X_4311_ _7414_/Q _4308_/S _4311_/A3 _4312_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor3_1
XFILLER_126_484 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_114_613 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_113_101 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5291_ _5624_/B _5759_/A1 _5431_/B _5292_/B _5291_/C _5293_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi221_1
Xoutput327 _7942_/Q wb_dat_o[24] VDD VSS gf180mcu_fd_sc_mcu7t5v0__buf_8
Xoutput338 _7501_/Q wb_dat_o[5] VDD VSS gf180mcu_fd_sc_mcu7t5v0__buf_8
XFILLER_99_357 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_7030_ _7133_/S _7030_/A2 _7030_/B _7933_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_4242_ _7732_/Q _6192_/A1 _4589_/A1 _7399_/Q _4243_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_68_700 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4173_ _7709_/Q _6141_/A1 hold119/I _7725_/Q _4174_/A4 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_7932_ _7932_/D _7961_/RN _7938_/CLK _7932_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_55_438 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_82_246 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_91_780 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7863_ _7863_/D _7901_/RN _7881_/CLK _7863_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffsnq_1
XFILLER_35_173 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_36_685 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7794_ _7794_/D _7901_/RN _7806_/CLK _7794_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
X_6814_ _7754_/Q _6644_/Z _6665_/Z _7746_/Q _6891_/C1 _7780_/Q _6815_/A4 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi222_1
XFILLER_23_357 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_50_121 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6745_ _7735_/Q _6830_/B _6889_/A2 _7703_/Q _6767_/C _6747_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi221_1
X_3957_ _7553_/Q _4284_/A1 _4427_/B _3958_/B2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_50_176 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_149_576 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3888_ _7781_/Q _6282_/A1 _6418_/A1 _7845_/Q _3892_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_6676_ _7700_/Q _6889_/A2 _6890_/A2 _7636_/Q _6677_/A4 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_5627_ _5741_/B _5627_/A2 _5627_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__and2_1
X_5558_ _5542_/Z _5557_/Z _5558_/B _5640_/B1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_105_602 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_172_590 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4509_ _4454_/Z _4521_/A2 _4509_/B hold704/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_5489_ _5548_/A1 _5150_/Z _5497_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_160_763 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_120_605 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7228_ _7228_/I0 _7948_/Q _7228_/S _7948_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_116_66 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7159_ _7159_/A1 _7159_/A2 _7159_/A3 _7159_/A4 _7160_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__or4_1
XFILLER_76_37 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_390 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_100_384 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_74_747 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_73_224 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2235 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2224 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2213 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2202 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_15_803 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_26_140 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_27_641 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2268 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2257 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2246 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1523 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1512 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1501 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_30 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_42_600 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_54_482 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2279 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_159_318 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_155_2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1567 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1556 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1545 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1534 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_41 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_25_63 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XPHY_52 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_63 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_74 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_1589 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1578 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_25_85 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_85 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_96 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_41_176 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_127_215 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_127_248 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_6_534 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_41_73 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_182_376 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_157_73 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_157_62 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_143_719 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_136_771 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_136_760 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_182_398 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_182_387 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_170_538 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_108_495 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_108_473 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_135_292 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_173_61 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_151_774 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_150_262 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_111_638 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_2_784 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_173_83 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_89_390 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_1_283 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_2_34 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_2_795 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_92_522 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_92_511 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_92_566 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_66_92 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_80_739 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_33_622 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_178_605 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_4860_ _4448_/Z _4862_/A2 _4860_/B _7523_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_3811_ _3801_/S hold629/Z _3811_/B _3843_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi21_4
XFILLER_60_463 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_60_474 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_32_165 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_177_148 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6530_ hold41/Z _6536_/A2 _6530_/B _7890_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_60_485 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_4791_ _7224_/I0 _7481_/Q _4795_/S _7481_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_118_204 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_70_2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3742_ _7346_/Q _7345_/Q _3751_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_2
X_3673_ hold66/Z _7273_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_6461_ hold380/Z _6468_/A2 _6462_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_173_376 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_161_505 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6392_ hold73/Z _6400_/A2 _6392_/B _7825_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_5412_ _5585_/A1 _5793_/A2 _5412_/B _5588_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_5343_ _5343_/A1 _5343_/A2 _5354_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_127_793 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_114_410 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_142_763 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_99_154 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xoutput168 _7982_/Z irq[0] VDD VSS gf180mcu_fd_sc_mcu7t5v0__buf_8
Xoutput179 _3695_/ZN mgmt_gpio_oeb[17] VDD VSS gf180mcu_fd_sc_mcu7t5v0__buf_8
XFILLER_102_605 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5274_ _5292_/B _5431_/B _5706_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_102_638 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7013_ _7896_/Q _7197_/A2 _6938_/I _7856_/Q _7014_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_68_530 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4225_ _7790_/Q _6316_/A1 _4604_/A1 _7405_/Q _4267_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_68_552 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4156_ _7767_/Q _6265_/A1 _5828_/A1 _7564_/Q _4604_/A1 _7406_/Q _4158_/A3 VDD VSS
+ gf180mcu_fd_sc_mcu7t5v0__aoi222_2
XFILLER_28_449 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_56_747 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4087_ _7848_/Q _6435_/A1 _6384_/A1 _7824_/Q _4090_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_36_460 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7915_ _7915_/D _7961_/RN _7940_/CLK _7915_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffsnq_2
X_7846_ _7846_/D _7901_/RN _7849_/CLK _7846_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffsnq_1
XFILLER_102_68 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_169_649 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_168_104 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_51_463 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4989_ _5006_/B _5006_/C _5344_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_4
X_7777_ _7777_/D _7901_/RN _7873_/CLK _7777_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_51_496 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6728_ _6728_/A1 _6728_/A2 _6728_/A3 _6728_/A4 _6728_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__and4_1
XFILLER_164_321 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_109_215 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6659_ _6878_/A2 _6665_/A2 _6659_/A3 _6659_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__and3_2
XFILLER_133_796 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_74_500 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_59_574 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_47_725 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2010 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2043 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2021 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2032 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_55_780 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2076 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2065 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2054 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1331 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1320 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_159_104 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2098 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2087 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1364 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1375 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1353 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1342 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_14_132 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_15_655 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_42_463 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1397 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1386 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_14_176 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_156_800 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_52_61 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xinput37 mgmt_gpio_in[10] input37/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
Xinput15 mask_rev_in[1] input15/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
Xinput26 mask_rev_in[2] input26/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_155_354 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xinput59 mgmt_gpio_in[30] input59/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
Xinput48 mgmt_gpio_in[20] input48/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_96_179 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4010_ _7720_/Q _6158_/A1 _6107_/A1 _7696_/Q _7680_/Q _6073_/A1 _4013_/A2 VDD VSS
+ gf180mcu_fd_sc_mcu7t5v0__aoi222_1
XFILLER_38_703 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_65_522 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_65_511 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_38_747 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_92_330 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_65_566 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5961_ hold527/Z _5970_/A2 _5962_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_18_460 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4912_ _4922_/A3 _4922_/A4 _4924_/A1 _4924_/A2 _4914_/A4 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand4_4
X_7700_ _7700_/D _7961_/RN _7701_/CLK _7700_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffsnq_1
X_7631_ _7631_/D _7901_/RN _7820_/CLK _7631_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
X_5892_ _4460_/Z _5902_/A2 _5892_/B _7590_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_61_783 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4843_ _4843_/A1 _7285_/A2 _4847_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_33_496 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_178_479 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_147_811 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7562_ _7562_/D input75/Z _7567_/CLK _7562_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
X_4774_ _4774_/A1 _7285_/A2 _4778_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_3725_ _5006_/C _5254_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_8
XFILLER_146_321 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6513_ hold41/Z _6519_/A2 _6513_/B _7882_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_20_179 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_7493_ _7493_/D _7912_/CLK _7493_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_6444_ hold334/Z _6451_/A2 _6445_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_119_557 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_146_398 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3656_ _7915_/Q _6905_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_2
XFILLER_161_357 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6375_ hold73/Z _6383_/A2 _6375_/B _7817_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_115_785 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5326_ _5326_/A1 _5326_/A2 _5326_/A3 _5326_/A4 _5354_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand4_1
XFILLER_142_582 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_5257_ _5394_/A1 _5005_/Z _5622_/A1 _5721_/C VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor3_1
XFILLER_130_744 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4208_ _7548_/Q _4427_/B _4284_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_180_29 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5188_ _5739_/A1 _5188_/A2 _5188_/A3 _5188_/A4 _5191_/B2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand4_1
XFILLER_29_747 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_29_769 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4139_ hold133/Z _4151_/A2 _4599_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_113_89 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_37_780 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_56_599 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_24_463 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7829_ _7829_/D _7901_/RN _7844_/CLK _7829_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_165_641 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_137_354 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_22_53 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_180_611 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_137_398 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_118_2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_106_763 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_78_102 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_121_766 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_121_799 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_93_105 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_78_179 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_19_224 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_90_812 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_170_95 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_74_385 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1150 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_15_430 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1183 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1172 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1161 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_15_496 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_30_400 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_43_783 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_179_93 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_147_107 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1194 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_128_321 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xhold618 _7825_/Q hold618/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
X_4490_ _4448_/Z _4504_/A2 _4490_/B _7355_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
Xhold607 _7536_/Q hold607/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
XFILLER_171_666 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_155_184 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_143_357 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xhold629 _3808_/Z hold629/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
XFILLER_170_176 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6160_ _4448_/Z _6174_/A2 _6160_/B _7716_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
XTAP_901 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_5111_ _5797_/B _5797_/C _5793_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_4
XFILLER_69_124 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_33_2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_912 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_923 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_934 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_6091_ hold625/Z _6106_/A2 _6092_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_945 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_956 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_967 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_978 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_5042_ _5548_/A1 _5043_/A2 _5042_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_97_499 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_84_105 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_989 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_81_812 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xclkbuf_leaf_51_csclk clkbuf_3_6__f_csclk/Z _7689_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_19_780 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6993_ _7831_/Q _7203_/A2 _7204_/B1 _7767_/Q _6997_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_179_733 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5944_ hold546/Z _5953_/A2 _5945_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_41_709 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5875_ _7583_/Q _5880_/A2 _5876_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_7614_ _7614_/D _7961_/RN _7707_/CLK _7614_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
X_4826_ _7226_/A1 _4828_/S _4826_/B _7500_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_138_129 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7545_ _7545_/D _7959_/RN _7545_/CLK _7545_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
Xclkbuf_leaf_66_csclk _7396_/CLK _7580_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_147_641 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_119_354 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_21_499 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4757_ hold617/Z _4758_/A2 _4758_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_146_173 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_146_151 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4688_ _3819_/Z _4448_/Z _4689_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_111_9 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7476_ _7476_/D _7961_/RN _7572_/CLK _7476_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
X_3708_ _7639_/Q _3708_/ZN VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_161_121 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_150_806 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6427_ hold391/Z _6434_/A2 _6428_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_3639_ _7414_/Q _4383_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_3
X_6358_ hold73/Z _6366_/A2 _6358_/B _7809_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_161_198 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5309_ _5309_/A1 _3723_/I _5344_/A1 _5433_/C _5495_/B2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand4_4
XFILLER_108_89 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_88_422 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_88_411 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6289_ hold530/Z _6298_/A2 _6290_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_102_232 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_48_308 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_130_596 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_124_33 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_88_488 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_84_37 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_90_108 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_72_812 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xclkbuf_leaf_19_csclk _7825_/CLK _7746_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_140_32 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_56_396 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_200 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_71_366 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_25_761 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_169_221 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_233 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_222 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_211 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_12_400 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_25_783 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_25_794 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_31_219 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_277 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_266 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_255 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_244 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_299 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_288 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_138_663 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_153_655 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_180_463 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_165_73 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_152_143 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_125_357 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_4_676 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_4_654 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_180_485 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_165_84 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xhold4 hold4/I hold4/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
XFILLER_121_596 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_79_499 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_47_330 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_63_812 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3990_ _3990_/A1 _3990_/A2 _3990_/A3 _3999_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor3_2
XFILLER_74_92 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_23_709 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_16_794 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5660_ _5079_/Z _5660_/A2 _5485_/B _5661_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor3_1
XFILLER_95_4 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_176_747 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_148_449 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_148_438 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_90_91 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_30_252 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4611_ _4448_/Z _4613_/A2 _4611_/B _7407_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_176_769 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5591_ _5474_/B _5591_/A2 _5454_/B _5656_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor3_1
XFILLER_129_641 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_117_803 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4542_ hold41/Z _4548_/A2 _4542_/B _7379_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_7330_ input75/Z _4334_/Z _7330_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__and2_1
X_7261_ _7261_/A1 _7261_/A2 _7262_/C VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
Xhold426 _7689_/Q hold426/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
Xhold415 _7735_/Q hold415/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
Xhold404 _7657_/Q hold404/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
X_4473_ hold453/Z _4487_/A1 hold454/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
Xhold437 _7746_/Q hold437/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
XFILLER_132_806 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_116_379 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6212_ hold728/Z _6225_/A2 _6213_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
Xhold459 _7568_/Q hold459/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
Xhold448 _7875_/Q hold448/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
XFILLER_171_496 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_143_176 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_131_349 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_7192_ _7192_/A1 _7192_/A2 _7192_/A3 _7209_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand3_1
X_6143_ _4448_/Z _6157_/A2 _6143_/B _7708_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_97_230 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_720 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_731 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_742 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_6074_ hold685/Z _6089_/A2 _6075_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_97_274 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_85_425 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_753 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_764 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_775 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_786 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_5025_ _5369_/B _5024_/Z _5535_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_100_747 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_85_447 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_797 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_72_108 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_93_491 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_81_631 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_54_29 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1919 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1908 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_6976_ _6976_/A1 _6976_/A2 _6976_/A3 _6976_/A4 _6977_/A4 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand4_1
XFILLER_26_569 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5927_ hold511/Z _5936_/A2 _5928_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_110_46 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5858_ hold41/Z _5868_/A2 _5858_/B _7575_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_182_717 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_166_257 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5789_ _5789_/A1 _5789_/A2 _5790_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_21_274 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4809_ _7228_/I0 _7492_/Q _4809_/S _7492_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_135_622 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_135_611 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_7528_ _7528_/D _7961_/RN _7625_/CLK _7528_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
X_7459_ _7459_/D _7901_/RN _7816_/CLK _7459_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_119_195 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_119_184 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_162_463 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_162_452 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_134_143 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_119_99 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_107_357 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_134_187 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_134_176 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_135_32 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_122_338 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_135_43 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_103_530 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_89_753 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_135_87 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_103_585 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_76_447 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_91_428 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_28_52 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_45_812 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_91_439 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_57_694 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_71_141 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_44_399 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_25_580 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_158_747 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_158_769 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_173_728 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_126_611 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_60_61 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_8_256 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_125_110 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_67_8 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_181_783 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_153_441 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_114_806 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_5_78 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_140_168 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_140_179 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_95_712 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_67_425 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_39_105 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_94_211 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_690 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_36_812 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_54_108 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_85_91 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6830_ _7739_/Q _6878_/A2 _6830_/B _6834_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_6761_ _7802_/Q _6883_/A2 _6883_/B1 _7786_/Q _6763_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_3973_ _7380_/Q hold114/I _6282_/A1 _7779_/Q _3985_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_5712_ _5104_/B _5669_/B _5712_/B _5716_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_149_736 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6692_ _6692_/A1 _6692_/A2 _6692_/A3 _6692_/A4 _6706_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand4_1
X_5643_ _5669_/B _5643_/A2 _5643_/B1 _5690_/A1 _5644_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_176_599 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_157_780 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_117_611 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5574_ _5705_/A2 _4996_/Z _5624_/A1 _5624_/B _5736_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_129_482 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xhold201 hold201/I _7654_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
X_7313_ input75/Z _4334_/Z _7313_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__and2_1
X_4525_ hold614/Z _4526_/A2 _4526_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
Xhold234 _7603_/Q hold234/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
XFILLER_144_463 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
Xhold212 _7734_/Q hold212/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
Xhold223 _7688_/Q hold223/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
X_7244_ _7518_/Q _7244_/A2 _7246_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
Xhold245 hold245/I _7848_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
Xhold278 _7634_/Q hold278/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
Xhold256 _7776_/Q hold256/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
Xhold267 hold267/I _7824_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
X_4456_ _4487_/A1 _4454_/Z _4456_/B hold737/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
Xhold289 _7852_/Q hold289/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
XFILLER_98_550 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4387_ _7448_/Q input89/Z _4387_/S _4387_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_7175_ _7476_/Q _7195_/A2 _7195_/B1 _7470_/Q _7195_/C1 _7383_/Q _7177_/A3 VDD VSS
+ gf180mcu_fd_sc_mcu7t5v0__aoi222_1
XFILLER_140_680 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_86_723 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_86_734 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_550 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_561 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_6126_ _4448_/Z _6140_/A2 _6126_/B _7700_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_100_544 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_86_756 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_58_458 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_572 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_583 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_594 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_100_555 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_100_566 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_39_650 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6057_ hold770/Z _6072_/A2 _6058_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_5008_ _5200_/B _5230_/A1 _5024_/A2 _5011_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor3_1
XFILLER_73_428 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1705 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_26_333 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_157_6 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1749 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1738 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1727 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1716 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_81_27 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_121_89 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_81_494 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6959_ _6959_/A1 _6959_/A2 _6959_/A3 _6959_/A4 _6977_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand4_1
XFILLER_53_185 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_182_558 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_5_237 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_5_215 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_182_569 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_107_132 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_163_783 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_135_496 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_123_636 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_100_2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_150_455 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_122_157 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_122_124 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_107_198 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_122_168 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_122_179 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_77_712 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_77_767 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_76_211 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_39_73 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_49_425 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_49_436 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_49_447 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_162_74 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_18_812 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_36_108 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_76_299 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_55_61 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_32_303 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_177_319 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_32_347 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xclkbuf_2_0__f_mgmt_gpio_in[4] clkbuf_0_mgmt_gpio_in[4]/Z _4418_/I1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_71_82 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_9_565 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_139_791 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_139_780 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_126_463 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xoutput306 _4424_/Z spimemio_flash_io0_di VDD VSS gf180mcu_fd_sc_mcu7t5v0__buf_8
Xoutput317 _7493_/Q wb_dat_o[15] VDD VSS gf180mcu_fd_sc_mcu7t5v0__buf_8
X_4310_ _7339_/Q _4294_/Z _4311_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_141_422 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5290_ _5687_/C _5350_/A3 _5290_/B _5291_/C VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi21_1
Xoutput328 _7943_/Q wb_dat_o[25] VDD VSS gf180mcu_fd_sc_mcu7t5v0__buf_8
XFILLER_5_760 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
Xoutput339 _7502_/Q wb_dat_o[6] VDD VSS gf180mcu_fd_sc_mcu7t5v0__buf_8
X_4241_ _7806_/Q _6350_/A1 _6124_/A1 _7700_/Q _4243_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_141_499 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4172_ _7717_/Q _6158_/A1 _4863_/A1 _7526_/Q _4174_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_7931_ _7931_/D _7961_/RN _7938_/CLK _7931_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_55_428 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_35_130 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_91_792 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7862_ _7862_/D _7901_/RN _7881_/CLK _7862_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffsnq_1
XFILLER_23_314 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_35_152 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_51_623 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7793_ _7793_/D _7901_/RN _7809_/CLK _7793_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
X_6813_ _7381_/Q _6882_/A2 _6894_/C1 _7836_/Q _6813_/C _6815_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi221_1
X_6744_ _7841_/Q _6894_/A2 _6659_/Z _7623_/Q _6747_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_3956_ _4206_/A1 _7228_/I0 _3958_/B1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_6675_ _7692_/Q _6881_/B1 _6882_/B1 _7652_/Q _6885_/B1 _7708_/Q _6677_/A3 VDD VSS
+ gf180mcu_fd_sc_mcu7t5v0__aoi222_1
XFILLER_149_566 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_109_408 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_5626_ _5391_/B _5706_/A2 _5626_/A3 _5625_/Z _5726_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand4_1
X_3887_ hold275/Z hold128/Z _6537_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_4
XFILLER_164_525 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_136_216 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_5557_ _5557_/A1 _5557_/A2 _5557_/A3 _5557_/A4 _5557_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__or4_1
XFILLER_129_290 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_117_430 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_145_783 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_144_260 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_117_496 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_117_485 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5488_ _5648_/A1 _5669_/B _5431_/B _5648_/B2 _5803_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_4508_ hold702/Z _4521_/A2 hold703/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_4439_ _7519_/Q _4338_/Z _7513_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_160_742 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7227_ _7227_/I0 _7947_/Q _7228_/S _7947_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_116_34 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_104_179 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_59_712 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7158_ _7158_/A1 _7158_/A2 _7158_/A3 _7158_/A4 _7159_/A4 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand4_1
XFILLER_86_531 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7089_ _7089_/A1 _7089_/A2 _7089_/A3 _7089_/A4 _7106_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand4_1
XFILLER_100_341 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6109_ _4448_/Z _6123_/A2 _6109_/B _7692_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
XTAP_391 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_380 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_132_33 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_86_586 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_74_737 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_18_108 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_46_439 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2225 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2214 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2203 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_39_491 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2269 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2258 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2247 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2236 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1524 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1513 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1502 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_92_37 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_20 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_31 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_25_20 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1557 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1546 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1535 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_42 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_25_53 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_53 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_64 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_148_2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1579 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1568 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_75 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_41_144 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XPHY_86 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_97 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_167_352 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_10_531 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_6_502 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_182_322 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_182_311 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_108_463 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_123_444 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_2_741 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_173_73 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_123_499 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_1_295 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_49_244 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_92_534 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_65_737 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_37_428 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_64_258 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_64_247 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_80_729 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_17_141 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_45_450 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_32_100 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3810_ hold23/Z _3808_/Z _3810_/S hold24/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_4790_ _7223_/A1 _4795_/S _4790_/B _7480_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_21_807 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3741_ _3734_/Z _3741_/A2 _3741_/B _7978_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_174_812 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3672_ hold45/Z _7268_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_173_333 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_6460_ hold73/Z _6468_/A2 _6460_/B _7857_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_6391_ hold618/Z _6400_/A2 _6392_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_5411_ _5669_/A1 _5793_/A2 _5292_/B _5482_/B2 _5411_/C _5413_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi221_1
XFILLER_63_2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_133_208 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_127_783 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5342_ _5621_/B _5724_/A2 _5759_/C _5721_/B _5343_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XFILLER_154_591 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_126_282 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_99_144 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_5273_ _5273_/A1 _5350_/A3 _5793_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_7012_ _7888_/Q _7196_/A2 _7196_/B1 _7638_/Q _7014_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_1
Xoutput169 _4432_/Z irq[1] VDD VSS gf180mcu_fd_sc_mcu7t5v0__buf_8
X_4224_ _7854_/Q _6452_/A1 _6333_/A1 _7798_/Q _4264_/A4 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_110_661 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_28_406 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4155_ hold275/Z _4155_/A2 _4527_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_110_672 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_83_523 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4086_ _7622_/Q _5954_/A1 _4231_/B1 input58/Z _4092_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_83_567 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7914_ _7914_/D _7961_/RN _7938_/CLK _7914_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_4
X_7845_ _7845_/D _7901_/RN _7901_/CLK _7845_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_23_144 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_7776_ _7776_/D _7901_/RN _7868_/CLK _7776_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffsnq_1
X_4988_ _5104_/B _5735_/A2 _5669_/A1 _5705_/A2 _4999_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_165_812 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3939_ _7812_/Q _6350_/A1 _5971_/A1 _7634_/Q _3940_/A4 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_6727_ _7800_/Q _6883_/A2 _6893_/B1 _7768_/Q _6891_/A2 _7824_/Q _6728_/A4 VDD VSS
+ gf180mcu_fd_sc_mcu7t5v0__aoi222_1
X_6658_ _6878_/A2 _6658_/A2 _6658_/A3 _6892_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor3_4
X_5609_ _5657_/A4 _5799_/A2 _5609_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_11_33 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_127_33 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6589_ _6590_/A1 _6665_/A2 _6830_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__and2_2
XFILLER_2_6 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_120_447 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_105_499 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_101_694 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_19_428 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_46_203 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2000 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_74_534 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_46_247 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2022 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2033 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2011 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2077 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2066 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2055 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2044 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1332 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1321 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1310 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_27_494 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2099 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2088 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1365 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1354 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1343 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1398 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1387 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1376 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_14_188 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_174_119 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_174_108 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_168_672 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_156_812 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_30_659 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_128_525 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_7_811 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
Xinput16 mask_rev_in[20] input16/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
Xinput27 mask_rev_in[30] input27/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
Xinput38 mgmt_gpio_in[11] input38/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
Xinput49 mgmt_gpio_in[21] input49/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_6_321 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_182_174 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_170_325 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_109_783 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_6_398 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_151_561 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_123_274 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_111_425 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_35_6 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_77_70 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_65_534 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_5960_ _4460_/Z _5970_/A2 _5960_/B hold186/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_4911_ _4924_/A3 _4924_/A4 _3727_/I _4914_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand3_2
X_5891_ hold196/Z _5902_/A2 _5892_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_178_414 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7630_ _7630_/D _7901_/RN _7797_/CLK _7630_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffsnq_2
X_4842_ _4376_/B _5520_/C _7279_/A2 _4842_/A4 _7506_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand4_1
XFILLER_60_250 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_21_615 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_33_486 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7561_ _7561_/D input75/Z _7561_/CLK _7561_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
X_4773_ _4454_/Z _4773_/A2 _4773_/B hold601/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_158_160 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3724_ _5006_/B _5394_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__inv_3
X_6512_ hold370/Z _6519_/A2 _6513_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_7492_ _7492_/D _7944_/CLK _7492_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_173_141 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6443_ hold73/Z _6451_/A2 _6443_/B _7849_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_107_709 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3655_ _7914_/Q _6908_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__inv_2
X_6374_ hold321/Z _6383_/A2 _6375_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_115_720 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_115_764 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_114_241 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5325_ _5624_/B _5624_/A2 _5724_/A2 _5685_/B _5326_/A4 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_88_615 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_519 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5256_ _5714_/B1 _5622_/A1 _5731_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_102_425 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_88_637 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_87_169 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4207_ _4207_/I0 _7549_/Q _4427_/B _7549_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_5187_ _5187_/A1 _5499_/A1 _5187_/A3 _5187_/A4 _5188_/A4 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor4_1
XFILLER_68_383 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_113_46 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_28_247 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_29_759 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4138_ _7741_/Q _6209_/A1 _4559_/A1 _7388_/Q _4158_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_56_534 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4069_ _4069_/A1 _4069_/A2 _7224_/I0 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_2
XFILLER_169_425 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_24_453 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7828_ _7828_/D _7901_/RN _7844_/CLK _7828_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_24_475 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_156_108 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_138_812 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7759_ _7759_/D _7901_/RN _7898_/CLK _7759_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffsnq_1
XFILLER_177_491 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_11_169 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_153_804 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_137_344 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_164_163 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_3_302 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_180_656 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_118_580 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_118_591 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_121_712 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_106_753 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_3_357 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_79_626 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_154_75 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_121_778 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_66_309 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_86_191 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_74_331 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_47_73 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_47_556 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_170_74 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_47_567 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_34_228 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1140 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1173 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1162 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1151 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_250 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_129_812 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1195 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1184 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_30_445 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_175_428 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_147_119 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_8_34 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_155_141 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_7_641 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xhold608 _7717_/Q hold608/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
Xhold619 _7587_/Q hold619/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
X_6090_ _6090_/A1 hold32/Z _6106_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_4
XFILLER_97_434 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_97_423 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5110_ _4996_/Z _5672_/A2 _5586_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_902 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_913 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_924 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_935 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_5041_ _5024_/Z _5041_/A2 _5533_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_112_756 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_946 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_957 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_968 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_97_478 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_26_2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_979 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_38_534 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xclkbuf_0_wb_clk_i wb_clk_i clkbuf_0_wb_clk_i/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_65_353 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_25_206 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_92_183 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_80_334 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6992_ _6992_/A1 _6992_/A2 _6992_/A3 _6992_/A4 _7001_/B1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand4_1
XFILLER_179_712 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_5943_ _4460_/Z _5953_/A2 _5943_/B hold152/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_5874_ _5874_/A1 hold32/Z _5880_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_2
XFILLER_80_389 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_61_570 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_138_108 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4825_ _7500_/Q _4828_/S _4826_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_7613_ _7613_/D _7961_/RN _7815_/CLK _7613_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_33_283 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_33_294 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_7544_ _7544_/D _7959_/RN _7545_/CLK _7544_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_146_130 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_119_344 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4756_ _4448_/Z _4758_/A2 _4756_/B _7466_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_146_163 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4687_ _7436_/Q _4718_/A1 _4690_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_3707_ _7647_/Q _3707_/ZN VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_7475_ _7475_/D _7961_/RN _7572_/CLK _7475_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
X_3638_ _7506_/Q _3810_/S VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_12
XFILLER_134_347 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6426_ hold73/Z _6434_/A2 _6426_/B _7841_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_161_144 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_6357_ hold503/Z _6366_/A2 _6358_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_5308_ _5498_/A2 _5687_/B _5510_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_103_712 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6288_ _4460_/Z _6298_/A2 _6288_/B _7776_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_130_531 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_349 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5239_ _5563_/B2 _5622_/A1 _5572_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_84_673 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_29_556 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_29_567 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_44_515 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_71_301 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_44_526 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_56_386 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_140_44 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_201 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_140_99 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_234 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_223 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_212 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_24_250 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_169_266 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XPHY_267 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_256 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_245 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_40_754 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_157_428 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_149_31 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_289 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_278 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_130_2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_33_64 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_149_64 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_8_449 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_137_141 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_165_494 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_152_155 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_98_209 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_67_618 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_66_117 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_58_72 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_181_73 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xhold5 hold5/I hold5/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
XFILLER_94_459 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_94_448 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_75_651 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_47_386 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_90_676 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_62_389 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_62_378 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_43_570 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_15_283 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4610_ hold664/Z _4613_/A2 _4611_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_175_247 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_175_236 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5590_ _5582_/Z _5590_/A2 _5590_/B _5639_/C VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_128_130 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_4541_ hold317/Z _4548_/A2 _4542_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_144_601 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_128_163 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7260_ _7520_/Q _7260_/A2 _7260_/B1 _7519_/Q _7261_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_143_111 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_116_314 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xhold416 _7687_/Q hold416/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
Xhold405 hold405/I _7657_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
X_4472_ _4487_/A1 hold41/Z _4472_/B hold491/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
Xhold427 _7876_/Q hold427/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
X_6211_ _4448_/Z _6225_/A2 _6211_/B _7740_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_143_144 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_32
Xhold449 _7780_/Q hold449/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
Xhold438 _7672_/Q hold438/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
X_7191_ _7510_/Q _7191_/A2 _7191_/B1 _7406_/Q _7192_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_6142_ hold638/Z _6157_/A2 _6143_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_710 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_112_531 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_721 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_732 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_743 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_6073_ _6073_/A1 hold32/Z _6089_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_4
XFILLER_97_286 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_754 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_765 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_776 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_5024_ _3728_/I _5024_/A2 _5024_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__xor2_1
XTAP_798 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_787 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_57_139 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_66_673 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_38_364 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_81_621 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_66_695 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_65_161 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_26_526 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_26_515 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1909 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_6975_ _7830_/Q _7203_/A2 _7204_/A2 _7838_/Q _6976_/A4 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_5926_ _4460_/Z _5936_/A2 _5926_/B hold150/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_139_428 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5857_ hold368/Z _5868_/A2 _5858_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_167_759 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_166_247 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5788_ _5412_/B _5788_/A2 _5789_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_21_286 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_22_798 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_4808_ _7227_/I0 _7491_/Q _4809_/S _7491_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_4739_ hold60/Z _4750_/I1 _4741_/S _7455_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_147_472 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_119_152 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_119_45 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_108_804 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_7527_ _7527_/D _7961_/RN _7625_/CLK _7527_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
X_7458_ _7458_/D _7901_/RN _7583_/CLK hold76/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
X_6409_ hold73/Z _6417_/A2 _6409_/B _7833_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_122_328 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_7389_ _7389_/D _7961_/RN _7874_/CLK _7389_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_1_636 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_146 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_76_459 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_178_2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_72_676 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_72_687 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_72_698 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_71_175 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_25_570 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_44_378 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_44_389 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_13_776 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_12_264 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_40_573 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_172_206 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_126_601 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_165_291 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_180_250 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_125_144 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_125_133 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_140_103 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
Xclkbuf_leaf_50_csclk clkbuf_3_6__f_csclk/Z _7673_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_4_463 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_79_231 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_121_361 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_79_286 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_39_139 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_36_802 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_75_470 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_48_684 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_48_673 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_47_194 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_6760_ _7842_/Q _6894_/A2 _6891_/A2 _7826_/Q _6763_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_35_378 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5711_ _5711_/A1 _5733_/A3 _5710_/Z _5717_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand3_1
X_3972_ _7360_/Q _4488_/A1 _6401_/A1 _7835_/Q _3996_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_93_2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6691_ _7759_/Q _6892_/A2 _6893_/C1 _7629_/Q _6692_/A4 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_176_534 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_148_247 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5642_ _5642_/A1 _5642_/A2 _5642_/A3 _5642_/A4 _5766_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand4_1
XFILLER_31_584 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_148_269 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5573_ _5573_/A1 _5759_/A1 _5573_/B _5573_/C _5732_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi211_1
Xhold202 _7694_/Q hold202/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
X_4524_ _4448_/Z _4526_/A2 _4524_/B _7371_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_7312_ input75/Z _4334_/Z _7312_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__and2_1
Xhold235 hold235/I _7603_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
Xhold213 hold213/I _6198_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
Xhold224 _7647_/Q hold224/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
X_7243_ _7243_/A1 _7277_/B _7243_/B _7950_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_171_283 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4455_ hold35/I hold2/Z hold3/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
Xhold268 _7811_/Q hold268/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
Xhold257 _7864_/Q hold257/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
Xhold246 _7349_/Q hold246/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
Xhold279 hold279/I _7634_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
X_4386_ _7449_/Q input91/Z _4387_/S _4386_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_7174_ _7523_/Q _7194_/A2 _7194_/B1 _7504_/Q _7194_/C1 _7409_/Q _7177_/A2 VDD VSS
+ gf180mcu_fd_sc_mcu7t5v0__aoi222_1
XFILLER_58_415 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_551 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_540 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_6125_ hold771/Z _6140_/A2 _6126_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_100_534 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_85_212 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_58_426 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_562 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_573 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_584 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_6056_ _6056_/A1 hold32/Z _6072_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_4
XFILLER_105_69 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_595 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_5007_ _4898_/Z _4915_/Z _5005_/Z _5151_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand3_2
XFILLER_66_481 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_38_161 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_121_35 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1706 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_26_345 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1739 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1728 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1717 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_81_473 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_14_529 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_54_676 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6958_ _7774_/Q _7200_/A2 _7189_/B1 _7684_/Q _7195_/B1 _7620_/Q _6959_/A4 VDD VSS
+ gf180mcu_fd_sc_mcu7t5v0__aoi222_1
XFILLER_179_361 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5909_ _4460_/Z hold276/I _5909_/B hold142/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_14_33 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_22_540 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6889_ _7526_/Q _6889_/A2 _6665_/Z _7538_/Q _6889_/C _6896_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi221_1
XFILLER_139_247 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_182_515 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_167_567 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_155_729 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_6_717 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_107_144 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_162_250 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_146_98 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_122_136 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_1_499 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_162_64 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_76_256 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_92_738 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_91_204 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_91_215 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_29_150 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_29_161 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_29_172 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_57_470 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_91_237 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_91_248 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_45_632 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_60_602 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_17_378 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_55_73 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_60_624 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_44_175 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_13_551 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_13_540 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_158_534 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_158_589 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_40_392 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xoutput307 _4425_/ZN spimemio_flash_io1_di VDD VSS gf180mcu_fd_sc_mcu7t5v0__buf_8
XFILLER_181_570 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xoutput329 _7944_/Q wb_dat_o[26] VDD VSS gf180mcu_fd_sc_mcu7t5v0__buf_8
XFILLER_5_783 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
Xoutput318 _7478_/Q wb_dat_o[16] VDD VSS gf180mcu_fd_sc_mcu7t5v0__buf_8
XFILLER_153_283 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4240_ _4240_/A1 _4240_/A2 _4240_/A3 _4240_/A4 _4283_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand4_2
X_4171_ _7522_/Q _4853_/A1 _4873_/A1 _7530_/Q _4174_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_95_532 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_67_212 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_82_204 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7930_ _7930_/D _7961_/RN _7940_/CLK _7930_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
X_7861_ _7861_/D _7901_/RN _7899_/CLK _7861_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
X_6812_ _6812_/A1 _6812_/A2 _6812_/A3 _6813_/C VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_36_676 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7792_ _7792_/D _7901_/RN _7806_/CLK _7792_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffsnq_1
XFILLER_90_281 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_50_101 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_50_112 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3955_ _3955_/A1 _3955_/A2 _3936_/Z _3955_/A4 _7228_/I0 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand4_4
X_6743_ _7615_/Q _6647_/Z _6887_/B1 _7679_/Q _6752_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_51_668 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6674_ _7782_/Q _6883_/B1 _6891_/C1 _7774_/Q _6674_/C _6677_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi221_1
XFILLER_176_353 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_136_206 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5625_ _5803_/A2 _5625_/A2 _5625_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__and2_1
X_3886_ _4153_/A1 _3886_/A2 _5988_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_4
X_5556_ _5642_/A4 _5649_/A4 _5557_/A4 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_144_250 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_132_412 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_132_401 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5487_ _5099_/B _5797_/A2 _5645_/A3 _5495_/B2 _5511_/C VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai22_1
X_4507_ _4448_/Z _4521_/A2 _4507_/B _7363_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_4438_ _5678_/A1 _4438_/A2 _7514_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_104_136 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_7226_ _7226_/A1 _7228_/S _7226_/B _7946_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_4369_ input97/Z input96/Z input99/Z input98/Z _4374_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor4_1
XFILLER_116_68 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7157_ _7765_/Q _7202_/C2 _7200_/B1 _7869_/Q _7158_/A4 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_98_392 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_7088_ _7713_/Q _7189_/A2 _7191_/B1 _7803_/Q _7089_/A4 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_86_543 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_6108_ hold624/Z _6123_/A2 _6109_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_59_779 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_392 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_370 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_381 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_6039_ _6039_/A1 hold32/Z _6055_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_4
XFILLER_74_727 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_73_215 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2226 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2215 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2204 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_132_67 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2259 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2248 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2237 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1514 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1503 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_21 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_10 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_15_805 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_42_602 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1547 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1536 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1525 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_14_337 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XPHY_32 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_43 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_54 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_65 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_41_112 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_54_484 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1569 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1558 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_76 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_87 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_98 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_22_370 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_155_515 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_10_521 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_22_392 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_182_301 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_127_228 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_127_217 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_41_53 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_163_570 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_157_86 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_135_283 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_123_423 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_96_307 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_173_63 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_96_329 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_49_212 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_92_513 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_73_771 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_18_676 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_45_495 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_177_106 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_20_318 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3740_ _4292_/B _3738_/Z _3741_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_119_707 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3671_ hold39/Z _7263_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_173_345 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6390_ _4460_/Z _6400_/A2 _6390_/B hold267/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_5410_ _5669_/A1 _5793_/A2 _5292_/B _5482_/B2 _5794_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_126_250 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5341_ _5645_/A3 _5495_/B2 _5721_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_114_412 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_56_2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_142_743 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_99_123 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5272_ _5199_/B _5201_/B _5338_/A1 _5369_/B _5350_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand4_4
X_7011_ _7646_/Q _7195_/A2 _7195_/B1 _7622_/Q _7188_/A2 _7377_/Q _7016_/A3 VDD VSS
+ gf180mcu_fd_sc_mcu7t5v0__aoi222_1
XFILLER_141_286 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_101_128 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4223_ _7838_/Q _6418_/A1 _4579_/A1 _7395_/Q _4256_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_4154_ hold275/Z _3881_/Z _5807_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_4085_ _7686_/Q _6090_/A1 _5828_/A1 _7565_/Q _6141_/A1 _7710_/Q _4092_/A2 VDD VSS
+ gf180mcu_fd_sc_mcu7t5v0__aoi222_2
XFILLER_83_513 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_55_215 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_56_727 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_83_546 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_83_557 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_83_535 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7913_ _7913_/D _7961_/RN _7938_/CLK _7913_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_4
XFILLER_102_37 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_102_26 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_24_602 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7844_ _7844_/D _7901_/RN _7844_/CLK _7844_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_24_646 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7775_ _7775_/D _7901_/RN _7897_/CLK _7775_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffsnq_1
XFILLER_51_432 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_51_443 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6726_ _7792_/Q _6893_/A2 _6892_/B1 _7726_/Q _6890_/B1 _7848_/Q _6728_/A3 VDD VSS
+ gf180mcu_fd_sc_mcu7t5v0__aoi222_1
X_4987_ _5669_/A1 _5705_/A2 _5706_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_3938_ input41/Z _5903_/A1 _6039_/A1 _7666_/Q _3940_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_3869_ _3869_/I _4653_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_6657_ _6878_/A2 _6661_/A3 _6658_/A3 _6893_/B1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor3_4
X_5608_ _5608_/A1 _5167_/B _5608_/B _5799_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_6588_ _7909_/Q _7908_/Q _6665_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_2
XFILLER_164_389 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5539_ _5543_/B _5153_/C _5539_/A3 _5552_/A4 _5546_/C VDD VSS gf180mcu_fd_sc_mcu7t5v0__or4_1
XFILLER_145_570 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_133_721 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_117_283 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_127_89 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_78_318 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7209_ _7210_/A2 _7209_/A2 _7209_/A3 _7209_/A4 _7210_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor4_1
XFILLER_101_651 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_59_565 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_86_384 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_59_576 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2001 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2023 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2034 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2012 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_160_2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2067 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2056 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2045 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1322 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1311 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1300 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_36_97 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_2089 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2078 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1366 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1355 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1344 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1333 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_30_605 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1399 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1388 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1377 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_498 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_168_651 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_128_504 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_128_515 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_10_340 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
Xinput17 mask_rev_in[21] input17/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
Xinput28 mask_rev_in[31] input28/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_182_142 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xinput39 mgmt_gpio_in[12] input39/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_108_250 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_123_286 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_97_638 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_96_148 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_77_384 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_37_215 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_92_321 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_53_708 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4910_ input97/Z input96/Z input99/Z input98/Z _4914_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand4_4
XFILLER_93_70 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5890_ _4454_/Z _5902_/A2 _5890_/B _7589_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_80_538 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_178_404 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4841_ _7506_/Q _7214_/A1 _4842_/A4 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_60_240 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_178_459 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_61_785 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_61_774 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_21_605 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_21_638 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7560_ _7560_/D input75/Z _7561_/CLK _7560_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffsnq_2
X_4772_ hold599/Z _4773_/A2 hold600/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_3723_ _3723_/I _5087_/C VDD VSS gf180mcu_fd_sc_mcu7t5v0__inv_4
XFILLER_174_621 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_158_183 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6511_ hold73/Z _6519_/A2 _6511_/B _7881_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_9_160 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_7491_ _7491_/D _7912_/CLK _7491_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_6442_ hold485/Z _6451_/A2 _6443_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_119_559 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3654_ _7911_/Q _6599_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_2
XFILLER_174_676 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_146_389 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_127_570 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6373_ _4460_/Z _6383_/A2 _6373_/B hold135/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_130_702 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5324_ _5624_/B _5624_/A2 _5647_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_88_605 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5255_ _5273_/A1 _5687_/C _5705_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_102_448 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4206_ _4206_/A1 _7221_/A1 _4206_/B _4207_/I0 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_57_19 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5186_ _5186_/A1 _5186_/A2 _5186_/A3 _5186_/A4 _5187_/A4 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand4_1
XFILLER_56_502 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_29_749 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4137_ hold133/Z _4217_/A2 _4559_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_113_69 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4068_ _4068_/A1 _4068_/A2 _4069_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_83_354 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_71_527 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_36_270 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_7827_ _7827_/D _7901_/RN _7851_/CLK _7827_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_12_605 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7758_ _7758_/D _7901_/RN _7826_/CLK _7758_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffsnq_1
X_7689_ _7689_/D _7961_/RN _7689_/CLK _7689_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
X_6709_ _7922_/Q _7133_/S _6710_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_22_11 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_165_632 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_138_33 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_164_175 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_138_66 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_106_743 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_98_37 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_133_540 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_105_231 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_120_212 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_105_286 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_79_638 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_160_392 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_93_107 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_74_321 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_19_215 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_170_64 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_74_365 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_35_708 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_47_96 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_28_782 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1141 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1130 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1174 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1163 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1152 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_63_84 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_63_73 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_30_402 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_42_262 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_43_785 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_179_73 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1196 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1185 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_11_682 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_156_676 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_128_389 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xhold609 _7528_/Q hold609/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
XFILLER_171_646 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_171_635 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_109_570 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_6_185 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_171_668 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_111_212 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_903 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_914 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_925 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_5040_ _5151_/A1 _5151_/A2 _5040_/B _5043_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi21_2
XFILLER_97_457 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_936 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_947 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_958 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_78_682 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_969 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_93_641 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_19_2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_38_524 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_6991_ _6991_/A1 _6991_/A2 _6992_/A4 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_92_173 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5942_ hold151/Z _5953_/A2 _5943_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_19_771 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5873_ _4448_/Z _5873_/A2 _5873_/B _7582_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_7612_ _7612_/D _7961_/RN _7815_/CLK _7612_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffsnq_1
XFILLER_61_593 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_61_582 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4824_ _7224_/I0 _7499_/Q _4828_/S _7499_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_159_481 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7543_ _7543_/D _7959_/RN _7545_/CLK hold23/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
X_4755_ hold696/Z _4758_/A2 _4756_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_3706_ _7655_/Q _3706_/ZN VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_174_451 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_162_602 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_146_153 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4686_ _4686_/A1 _5903_/A2 _4686_/B1 _3819_/Z hold12/Z _4718_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi221_4
X_7474_ _7474_/D _7961_/RN _7572_/CLK _7474_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_162_646 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6425_ hold365/Z _6434_/A2 _6426_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_3637_ _7344_/Q _3744_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__inv_1
X_6356_ _4460_/Z _6366_/A2 _6356_/B _7808_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_5307_ _5307_/A1 _5307_/A2 _5650_/A3 _5433_/C _5307_/B2 _5356_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai32_1
XFILLER_103_724 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_68_29 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_317 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_142_392 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6287_ hold256/Z _6298_/A2 _6288_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_5238_ _5200_/B _3727_/I _5421_/A1 _5433_/C _5622_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand4_4
XFILLER_124_46 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5169_ _5643_/A2 _5672_/A2 _5793_/A2 _5167_/B _5171_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_84_28 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_69_682 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_56_321 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_140_34 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_84_685 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_17_33 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_83_195 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_71_357 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_17_77 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_169_212 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_224 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_213 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_202 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_12_402 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_268 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_257 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_246 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_235 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_33_32 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_40_744 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_169_278 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_279 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_137_131 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_123_2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_138_676 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_4_601 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_152_112 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_152_101 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_3_100 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_152_134 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_106_540 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_3_144 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_140_329 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_140_318 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_121_565 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_48_811 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
Xhold6 hold6/I hold6/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
XFILLER_66_129 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_47_321 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_75_641 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_47_354 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_74_162 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_74_195 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_50_519 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_15_295 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_175_215 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4540_ hold73/Z _4548_/A2 _4540_/B _7378_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_128_153 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
Xhold417 _7673_/Q hold417/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
Xhold406 _7705_/Q hold406/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
X_4471_ hold489/Z _4487_/A1 hold490/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_6210_ hold652/Z _6225_/A2 _6211_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
Xhold439 hold439/I _7672_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
Xhold428 _7617_/Q hold428/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
X_7190_ _7402_/Q _7190_/A2 _7190_/B1 _7469_/Q _7190_/C1 _7526_/Q _7192_/A2 VDD VSS
+ gf180mcu_fd_sc_mcu7t5v0__aoi222_1
X_6141_ _6141_/A1 hold32/Z _6157_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_4
XFILLER_131_307 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_124_370 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_98_733 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_700 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_124_392 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_98_744 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_711 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_722 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_733 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_6072_ hold90/Z _6072_/A2 _6072_/B hold345/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_98_788 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_744 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_755 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_766 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_777 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_5023_ _5338_/A1 _5024_/A2 _5040_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_100_738 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_799 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_788 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_38_321 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_38_376 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6974_ _7644_/Q _7195_/A2 _7190_/B1 _7612_/Q _6976_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_53_346 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_53_357 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5925_ hold148/Z _5936_/A2 hold149/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_80_176 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_110_37 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5856_ hold26/Z hold32/Z _5868_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_4
XFILLER_167_716 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4807_ _4807_/A1 _4809_/S _4807_/B _7490_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_5787_ _5787_/A1 _5787_/A2 _5787_/A3 _7544_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand3_1
X_4738_ hold63/Z _4749_/I1 _4741_/S _7454_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_7526_ _7526_/D _7961_/RN _7650_/CLK _7526_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_174_281 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4669_ _4685_/A1 hold74/Z _4669_/B hold75/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_7457_ _7457_/D _7901_/RN _7816_/CLK _7457_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_150_605 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_134_156 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6408_ hold538/Z _6417_/A2 _6409_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_122_318 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7388_ _7388_/D _7961_/RN _7531_/CLK _7388_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_150_649 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_6339_ _4460_/Z _6349_/A2 _6339_/B hold264/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_103_532 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_135_67 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_8009_ _8009_/I _8009_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_88_287 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_28_54 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_28_65 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_29_354 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_57_641 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_151_88 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_56_195 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_13_700 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_44_53 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_44_368 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_44_64 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_157_215 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_157_248 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_13_799 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_8_247 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_153_432 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_126_668 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_181_785 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_141_638 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_141_627 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_180_295 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_106_392 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_95_703 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_94_202 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_95_769 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_10_6 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_47_140 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_85_93 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3971_ _7899_/Q _6537_/A1 hold108/I _8009_/I _3998_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_90_463 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_16_560 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_35_357 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_35_368 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_5710_ _5710_/A1 _5710_/A2 _5710_/A3 _5710_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__and3_1
XFILLER_149_705 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_62_176 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6690_ _7823_/Q _6891_/A2 _6891_/B1 _7669_/Q _6892_/B1 _7725_/Q _6692_/A3 VDD VSS
+ gf180mcu_fd_sc_mcu7t5v0__aoi222_1
X_5641_ _5641_/A1 _5641_/A2 _5558_/B _5747_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_86_2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_31_574 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_157_771 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5572_ _4996_/Z _5608_/B _5572_/B _5572_/C _5716_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi211_2
XFILLER_129_495 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4523_ hold701/Z _4526_/A2 _4524_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_7311_ input75/Z _4334_/Z _7311_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__and2_1
X_7242_ _7242_/A1 _7280_/A2 _7277_/B _7242_/C _7243_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi211_1
Xhold214 hold214/I _7734_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
Xhold203 hold203/I _7694_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
Xhold225 hold225/I _6013_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
XFILLER_172_796 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_4454_ hold35/Z hold2/Z _4454_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__and2_4
Xhold269 _7745_/Q hold269/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
Xhold236 _7821_/Q hold236/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
XFILLER_132_605 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xhold258 hold258/I _7864_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
XFILLER_116_189 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_104_329 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_104_318 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xhold247 hold247/I _4462_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
X_4385_ _5678_/A1 _4338_/Z _7215_/C _7516_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_7173_ _7395_/Q _7193_/A2 _7193_/B1 _7472_/Q _7193_/C1 _7531_/Q _7177_/A1 VDD VSS
+ gf180mcu_fd_sc_mcu7t5v0__aoi222_1
X_6124_ _6124_/A1 hold32/Z _6140_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_4
XTAP_530 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_541 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_552 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_6055_ hold90/Z _6055_/A2 _6055_/B hold220/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_86_747 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_563 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_574 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_585 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_5006_ _3722_/I _3723_/I _5006_/B _5006_/C _5024_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai211_4
XTAP_596 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_27_803 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_39_641 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_66_460 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_39_685 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_54_600 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_66_493 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_1729 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1718 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1707 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_6957_ _7814_/Q _7207_/A2 _7190_/C1 _7700_/Q _6959_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_54_666 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_81_496 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_41_349 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_139_215 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5908_ hold140/Z hold276/I hold141/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_6888_ _6888_/A1 _6888_/A2 _6888_/A3 _6888_/A4 _6888_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__and4_1
X_5839_ hold459/Z _5840_/A2 _5840_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_155_719 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_108_602 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_10_747 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_182_527 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7509_ _7509_/D _7961_/RN _7510_/CLK _7509_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_30_33 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_30_55 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_163_785 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_146_33 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_123_638 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_122_104 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_146_77 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xhold770 _7668_/Q hold770/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
XFILLER_122_159 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_89_574 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_77_703 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_131_682 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_130_192 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_85_780 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_57_482 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_72_463 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_17_357 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_17_368 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_44_143 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_32_316 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_32_327 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_71_73 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_9_512 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_9_567 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xoutput308 _8008_/Z spimemio_flash_io2_di VDD VSS gf180mcu_fd_sc_mcu7t5v0__buf_8
XFILLER_114_605 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_99_316 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_4_250 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xoutput319 _7479_/Q wb_dat_o[17] VDD VSS gf180mcu_fd_sc_mcu7t5v0__buf_8
XFILLER_114_649 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4170_ _4167_/Z _4170_/A2 _4170_/A3 _4204_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand3_2
XFILLER_68_747 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_96_81 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_68_769 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_68_758 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_83_728 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_48_460 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7860_ _7860_/D _7901_/RN _7901_/CLK _7860_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_76_791 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_6811_ _7666_/Q _6885_/A2 _6893_/B1 _7772_/Q _6812_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_91_783 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_91_772 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_91_761 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_90_271 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_90_260 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7791_ _7791_/D _7961_/RN _7791_/CLK _7791_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffsnq_1
XFILLER_63_496 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_51_625 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3954_ _3954_/A1 _3954_/A2 _3954_/A3 _3954_/A4 _3955_/A4 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor4_4
X_6742_ _6742_/A1 _6742_/A2 _6742_/A3 _6753_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_50_157 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_176_321 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_149_546 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_3885_ hold128/Z hold133/Z _6401_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_4
X_6673_ _6673_/A1 _6673_/A2 _6673_/A3 _6674_/C VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_50_179 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_5624_ _5624_/A1 _5624_/A2 _5648_/B2 _5624_/B _5626_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai31_1
X_5555_ _5179_/B _5793_/A2 _5555_/B _5555_/C _5649_/A4 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XFILLER_172_582 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_5486_ _5543_/B _5504_/B1 _5553_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_145_785 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_144_262 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_117_465 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4506_ hold763/Z _4521_/A2 _4507_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_4437_ _7518_/Q _4338_/Z _7515_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_160_744 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_105_638 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7225_ _7946_/Q _7228_/S _7226_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_101_800 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_7156_ _7805_/Q _7191_/B1 _7188_/A2 _7382_/Q _7158_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_4368_ _4368_/A1 _4368_/A2 _4368_/A3 _4372_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor3_1
XFILLER_76_29 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6107_ _6107_/A1 hold32/Z _6123_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_4
X_4299_ _7343_/Q _4383_/A1 _4297_/Z _4300_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand3_1
X_7087_ _7689_/Q _7189_/B1 _7189_/C1 _7657_/Q _7089_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_100_343 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_100_321 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_393 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_371 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_382 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_6038_ hold90/Z _6038_/A2 _6038_/B hold339/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_74_717 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_67_780 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2216 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2205 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_67_791 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2249 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2238 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2227 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_162_6 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_132_79 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_1515 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1504 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_22 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_11 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_54_463 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7989_ _7989_/I _7989_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_1548 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1537 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1526 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_33 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_44 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_26_176 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_26_198 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XPHY_55 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_41_102 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_42_636 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_54_474 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_168_800 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1559 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_66 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_77 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_88 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_179_181 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_99 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_167_354 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_182_324 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xclkbuf_leaf_64_csclk _7961_/CLK _7701_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_182_368 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_163_560 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_151_766 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_151_799 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_110_118 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_104_693 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_1_286 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_49_224 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_106_80 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_77_544 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_2_37 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_77_588 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_65_739 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_18_666 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
Xclkbuf_leaf_17_csclk _7592_/CLK _7889_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_73_783 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_158_321 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_82_94 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_32_179 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3670_ hold71/Z _7258_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_158_398 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_173_357 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_161_519 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5340_ _5689_/A2 _5687_/B _5504_/A3 _5618_/B1 _5498_/A2 _5759_/C VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai32_1
X_5271_ _3728_/I _5022_/B _5271_/A3 _5431_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor3_4
XFILLER_5_570 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_49_2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_102_619 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_7010_ _7694_/Q _7194_/A2 _7194_/B1 _7662_/Q _7194_/C1 _7808_/Q _7016_/A2 VDD VSS
+ gf180mcu_fd_sc_mcu7t5v0__aoi222_1
XFILLER_88_809 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4222_ _7774_/Q _6282_/A1 _4584_/A1 _7397_/Q _4264_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_68_500 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4153_ _4153_/A1 hold107/Z _4812_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_4084_ _4084_/A1 _4084_/A2 _4084_/A3 _4084_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__and3_1
XFILLER_28_408 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_49_780 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7912_ _7912_/D _7961_/RN _7912_/CLK _7912_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffsnq_4
XFILLER_71_709 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_36_463 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7843_ _7843_/D _7901_/RN _7873_/CLK _7843_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_63_271 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_4986_ _4993_/B _5647_/A2 _5705_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_4
X_7774_ _7774_/D _7901_/RN _7898_/CLK _7774_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffsnq_1
X_6725_ _7808_/Q _6880_/B1 _6665_/Z _7742_/Q _6728_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_3937_ _7780_/Q _6282_/A1 _6248_/A1 _7764_/Q _6401_/A1 _7836_/Q _3940_/A2 VDD VSS
+ gf180mcu_fd_sc_mcu7t5v0__aoi222_2
XFILLER_51_499 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_177_641 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_149_354 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_176_162 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3868_ hold123/Z _3925_/A2 hold127/Z _3963_/A4 _3869_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__or4_4
X_6656_ _6878_/A2 _6664_/A3 _6658_/A3 _6891_/C1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor3_4
X_3799_ _7341_/Q _7414_/Q _3799_/B hold131/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi21_2
X_5607_ _5648_/A2 _5606_/B _5657_/A4 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_6587_ _6636_/A1 _6587_/A2 _6587_/B _7909_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_5538_ _5538_/A1 _5548_/A1 _5643_/B1 _5150_/Z _5652_/A4 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand4_1
XFILLER_133_700 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_11_35 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_160_530 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_127_46 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_127_35 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_118_796 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_133_777 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5469_ _5735_/A2 _5643_/A2 _5672_/A2 _4996_/Z _5749_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_7208_ _7208_/A1 _7208_/A2 _7208_/A3 _7208_/A4 _7209_/A4 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand4_1
XFILLER_160_585 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_59_522 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_59_511 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7139_ _7821_/Q _7207_/A2 _7201_/A2 _7755_/Q _7140_/A4 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_101_641 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_59_555 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2024 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2013 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2002 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_27_430 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_36_54 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2068 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2057 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2046 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2035 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1323 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1312 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1301 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_27_496 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_55_783 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2079 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_153_2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1356 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1345 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1334 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_82_591 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_14_124 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_15_647 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_159_118 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1389 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1367 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1378 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_14_179 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_52_53 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_167_162 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_155_302 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
Xinput18 mask_rev_in[22] input18/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_155_357 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xinput29 mask_rev_in[3] input29/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_6_378 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_124_744 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_123_221 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_123_210 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_6_389 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_124_755 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_123_232 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_96_105 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_93_812 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_18_463 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4840_ _7517_/D _7513_/Q _7515_/Q _7514_/Q _7279_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor4_2
XFILLER_45_282 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_178_449 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_61_797 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_20_105 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_159_641 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_147_803 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1890 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_6510_ hold372/Z _6519_/A2 _6511_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_4771_ _4448_/Z _4773_/A2 _4771_/B _7472_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_33_499 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3722_ _3722_/I _5309_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_8
X_7490_ _7490_/D _7944_/CLK _7490_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_158_195 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_6441_ _4460_/Z _6451_/A2 _6441_/B hold245/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_146_346 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_119_538 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3653_ _7434_/Q _4352_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_2
X_6372_ _7816_/Q _6383_/A2 _6373_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_5323_ _5724_/B _5648_/B2 _5724_/A2 _5624_/B _5326_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_5254_ _5006_/B _5254_/A2 _5254_/A3 _5433_/C _5409_/B2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand4_4
XFILLER_87_105 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_130_747 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5185_ _5666_/A1 _5669_/B _5185_/B _5512_/B _5186_/A4 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi211_1
X_4205_ _7548_/Q _4206_/A1 _4206_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_110_460 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_84_812 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_3_80 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4136_ hold113/Z _4155_/A2 _6243_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_4067_ _4067_/A1 _4067_/A2 _4067_/A3 _4067_/A4 _4068_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand4_1
XFILLER_37_783 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7826_ _7826_/D _7901_/RN _7826_/CLK _7826_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_52_742 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4969_ _5774_/A1 _5709_/A1 _4969_/B _4969_/C _4999_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai211_1
X_7757_ _7757_/D _7961_/RN _7874_/CLK _7757_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_149_140 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7688_ _7688_/D _7961_/RN _7692_/CLK _7688_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
X_6708_ _7433_/Q _7921_/Q _6708_/B _6710_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_149_184 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_22_45 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6639_ _6878_/A2 _6663_/A4 _6658_/A3 _6883_/B1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor3_4
XFILLER_137_357 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_125_508 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_133_563 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_160_382 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_101_460 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_93_119 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_87_661 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_75_812 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_59_374 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_19_238 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1120 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1131 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1164 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1153 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1142 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1197 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1186 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1175 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_15_488 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_15_499 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_42_274 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_175_419 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_156_600 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_7_632 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_10_193 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_171_658 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_170_179 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_97_425 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_904 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_915 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_926 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_112_747 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_111_246 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_2_392 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_937 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_948 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_959 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_84_108 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_66_812 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_65_311 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_93_653 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6990_ _6990_/A1 _6990_/A2 _6990_/A3 _6990_/A4 _6991_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand4_1
XFILLER_38_569 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5941_ _4454_/Z _5953_/A2 _5941_/B _7613_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_19_783 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_179_725 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_178_213 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5872_ hold558/Z _5873_/A2 _5873_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_178_257 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7611_ _7611_/D _7961_/RN _7694_/CLK _7611_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_21_425 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4823_ _7223_/A1 _4828_/S _4823_/B _7498_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_7542_ _7542_/D _7959_/RN _7545_/CLK hold18/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
X_4754_ _4754_/A1 _7285_/A2 _4758_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_3705_ _7663_/Q _3705_/ZN VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_7473_ _7473_/D _7961_/RN _7510_/CLK _7473_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_174_463 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_146_132 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4685_ _4685_/A1 _4685_/A2 hold98/Z hold99/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_119_357 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6424_ _4460_/Z _6434_/A2 _6424_/B _7840_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_3636_ _7553_/Q _4002_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_162_669 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6355_ hold136/Z _6366_/A2 _6356_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_108_37 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5306_ _5645_/A1 _5421_/B1 _5650_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_115_585 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6286_ _4454_/Z _6298_/A2 _6286_/B _7775_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_5237_ _5433_/C _5621_/B _5237_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_88_447 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_102_246 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_29_503 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_57_812 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5168_ _5643_/A2 _5672_/A2 _5673_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_5099_ _4993_/C _5663_/A1 _5099_/B _5573_/C VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_17_709 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4119_ hold113/Z _4217_/A2 _4604_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_140_46 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_225 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_214 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_203 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_24_263 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_52_572 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7809_ _7809_/D _7901_/RN _7809_/CLK _7809_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XPHY_258 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_247 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_236 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_157_408 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_138_600 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_269 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_165_496 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_153_647 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_137_176 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_125_327 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_116_2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_4_646 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_165_98 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_152_179 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_79_425 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_3_156 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_133_382 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_66_108 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xhold7 hold7/I hold7/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
XFILLER_114_91 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_47_377 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_74_84 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_16_742 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_31_712 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_50_509 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_130_90 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_30_211 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_156_463 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4470_ hold41/Z _4749_/I1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_128_176 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xhold407 _7829_/Q hold407/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
Xhold418 hold418/I _7673_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
XFILLER_143_135 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xhold429 hold429/I _7617_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
XFILLER_99_81 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_171_499 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6140_ hold90/Z _6140_/A2 _6140_/B _7707_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
XTAP_701 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_152_691 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_124_382 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_112_544 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_712 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_31_2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_723 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_734 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_6071_ hold344/Z _6072_/A2 _6072_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_112_555 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_112_566 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_745 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_756 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_767 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_39_812 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5022_ _5338_/A1 _5024_/A2 _5022_/B _5151_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_2
XFILLER_85_428 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_778 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_38_311 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_789 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_65_141 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_66_686 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_65_152 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_26_517 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_81_645 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6973_ _7708_/Q _7189_/A2 _7193_/B1 _7628_/Q _6938_/I _7854_/Q _6976_/A2 VDD VSS
+ gf180mcu_fd_sc_mcu7t5v0__aoi222_1
X_5924_ _4454_/Z _5936_/A2 _5924_/B _7605_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_179_566 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5855_ _5855_/A1 _4448_/Z _5855_/B hold12/Z hold13/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XFILLER_22_734 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4806_ _7490_/Q _4809_/S _4807_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_5786_ _7544_/Q _5520_/C _5786_/B1 _5792_/B1 _5786_/C1 _5802_/A1 _5787_/A3 VDD VSS
+ gf180mcu_fd_sc_mcu7t5v0__aoi222_1
XFILLER_182_709 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4737_ hold82/Z _4748_/I1 _4741_/S _7453_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_7525_ _7525_/D _7961_/RN _7650_/CLK _7525_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_175_783 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_174_271 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7456_ _7456_/D _7901_/RN _7743_/CLK _7456_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_162_400 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4668_ _7461_/Q hold55/Z _4668_/B hold74/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_147_496 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_119_176 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_119_69 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6407_ _4460_/Z _6417_/A2 _6407_/B _7832_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_102_8 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_134_168 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_134_179 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_89_712 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7387_ _7387_/D _7961_/RN _7510_/CLK _7387_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
X_4599_ _4599_/A1 _7285_/A2 _4603_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_6338_ hold263/Z _6349_/A2 _6339_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_104 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_1_638 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_95_39 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_95_28 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_89_778 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6269_ _4454_/Z _6281_/A2 _6269_/B _7767_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_48_108 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_130_385 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_130_396 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8008_ _8008_/I _8008_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_88_299 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_48_119 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_69_491 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_28_44 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_28_33 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_84_483 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_84_450 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_72_601 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_71_122 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_44_325 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_72_678 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_71_144 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_25_561 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_71_177 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_13_712 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_25_594 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_158_717 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_40_531 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_157_227 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_40_575 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_173_709 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_138_463 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_60_53 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_125_102 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_180_241 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_180_230 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_126_658 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_99_509 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_140_105 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_180_285 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_153_499 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_69_73 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_121_363 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_95_759 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_79_288 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_67_428 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_682 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_39_119 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_94_247 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_47_130 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3970_ input49/Z _4275_/A2 _5886_/A1 input57/Z _4239_/A2 input25/Z _3998_/A2 VDD
+ VSS gf180mcu_fd_sc_mcu7t5v0__aoi222_1
XFILLER_90_475 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_16_550 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_62_188 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_176_547 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_5640_ _5640_/A1 _5520_/C _5640_/B1 _5640_/B2 _7541_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_5571_ _5585_/A1 _5658_/B _5585_/B _5585_/C _5784_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XFILLER_79_2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_157_783 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_8_771 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7310_ input75/Z _4334_/Z _7310_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__and2_1
X_4522_ _4522_/A1 _7285_/A2 _4526_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_7241_ _7241_/A1 _7241_/A2 _7242_/C VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_4453_ hold1/Z _3810_/S hold2/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_156_282 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
Xhold204 _7715_/Q hold204/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
Xhold215 _7678_/Q hold215/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
Xhold226 hold226/I _7647_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
Xhold259 _7820_/Q hold259/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
Xhold237 _7683_/Q hold237/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
XFILLER_116_179 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xhold248 hold248/I _7349_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
X_4384_ _7511_/Q _7214_/A2 _7215_/C VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_171_296 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_98_531 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7172_ _7172_/A1 _7172_/A2 _7172_/A3 _7178_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand3_1
X_6123_ hold90/Z _6123_/A2 _6123_/B _7699_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
XTAP_531 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_520 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_542 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_6054_ hold218/Z _6055_/A2 hold219/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_140_672 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_553 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_564 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_575 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_5005_ _3722_/I _3723_/I _5005_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__or2_2
XTAP_586 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_597 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_93_280 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_66_483 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_38_196 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_53_122 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_1719 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1708 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_81_475 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6956_ _7676_/Q _7191_/A2 _7204_/B1 _7766_/Q _6959_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_53_144 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5907_ _4454_/Z hold276/Z _5907_/B _7597_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_34_380 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6887_ _7469_/Q _6647_/Z _6887_/B1 _7510_/Q _6887_/C _6888_/A4 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi221_1
XFILLER_139_227 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5838_ hold41/Z _5840_/A2 _5838_/B _7567_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_155_709 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5769_ _5769_/A1 _5769_/A2 _5651_/Z _5769_/A4 _5770_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__and4_1
XFILLER_22_597 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_7508_ _7508_/D _7961_/RN _7531_/CLK _7508_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_162_252 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_146_45 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_135_488 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7439_ _7439_/D _7961_/RN _7673_/CLK _7988_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_146_89 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
Xhold760 _7846_/Q hold760/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
XFILLER_135_499 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
Xhold771 _7700_/Q hold771/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
XFILLER_89_542 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_49_428 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_76_258 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_76_247 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_29_141 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_17_336 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_44_100 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_44_188 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_158_514 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_111_70 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_13_542 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_13_586 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_139_783 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_154_764 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
Xoutput309 _8009_/Z spimemio_flash_io3_di VDD VSS gf180mcu_fd_sc_mcu7t5v0__buf_8
XFILLER_5_785 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_4_262 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_110_812 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_95_567 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_95_578 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_63_420 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_48_494 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6810_ _7804_/Q _6883_/A2 _6883_/B1 _7788_/Q _6812_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_90_250 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_35_144 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_90_283 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7790_ _7790_/D _7901_/RN _7834_/CLK _7790_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffsnq_1
XFILLER_35_177 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_177_812 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3953_ _3953_/A1 _3953_/A2 _3953_/A3 _3953_/A4 _3954_/A4 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand4_2
X_6741_ _7378_/Q _6882_/A2 _6880_/A2 _7817_/Q _6742_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_149_536 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3884_ hold146/Z hold133/Z _6418_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_4
X_6672_ _7790_/Q _6893_/A2 _6659_/Z _7620_/Q _6673_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_31_361 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5623_ _5623_/A1 _5620_/B _5790_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_5554_ _5641_/A1 _5641_/A2 _5652_/A4 _5769_/A2 _5557_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand4_1
XFILLER_117_422 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5485_ _5680_/A1 _5779_/B1 _5485_/B _5504_/B1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_4505_ _4505_/A1 _7285_/A2 _4521_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_4
XFILLER_160_734 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_117_499 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7224_ _7224_/I0 _7945_/Q _7228_/S _7945_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_4436_ _7979_/Q input75/Z _4436_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__or2_1
X_4367_ _4367_/A1 _4367_/A2 _4367_/A3 _4372_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor3_1
XFILLER_132_469 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_116_37 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_7155_ _7901_/Q _7197_/A2 _7195_/B1 _7627_/Q _7158_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_113_694 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6106_ hold90/Z _6106_/A2 _6106_/B _7691_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_101_812 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4298_ _7343_/Q _4309_/S _4301_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_7086_ _7681_/Q _7191_/A2 _7190_/B1 _7617_/Q _7190_/A2 _7795_/Q _7089_/A2 VDD VSS
+ gf180mcu_fd_sc_mcu7t5v0__aoi222_1
XFILLER_86_567 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_86_534 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_58_247 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_372 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_394 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_383 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_6037_ hold338/Z _6038_/A2 _6038_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_73_206 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2217 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2206 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_100_388 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2239 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2228 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1505 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_92_29 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_12 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_54_453 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_7988_ _7988_/I _7988_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_1538 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1527 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1516 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_81_283 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_23 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_34 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_45 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_26_188 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_56 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_1549 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_67 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_78 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_41_136 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6939_ _6953_/A2 _6950_/A2 _6941_/A2 _7193_/C1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor3_4
XPHY_89 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_10_534 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_41_22 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_157_44 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_163_550 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_151_712 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xclkbuf_0_csclk _4416_/ZN clkbuf_0_csclk/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_151_723 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_150_211 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_123_425 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_9_2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_2_733 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_151_778 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
Xhold590 _7522_/Q hold590/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
XFILLER_110_108 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_77_523 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_2_788 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_18_623 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_17_144 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_72_250 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_33_626 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_60_456 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_60_467 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_119_709 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_158_388 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_146_528 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_9_354 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5270_ _5292_/B _5624_/B _5391_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_102_609 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4221_ _7355_/Q _4488_/A1 _4554_/A1 _7385_/Q _4264_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_68_534 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4152_ hold275/Z hold156/Z _4549_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_4083_ _7718_/Q _6158_/A1 _4083_/B _4084_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_7911_ _7911_/D _7961_/RN _7912_/CLK _7911_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffsnq_4
XFILLER_91_570 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7842_ _7842_/D _7901_/RN _7897_/CLK _7842_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_168_108 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_4985_ _5022_/B _4943_/Z _5647_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_4
X_7773_ _7773_/D _7901_/RN _7877_/CLK _7773_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_63_283 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6724_ _7662_/Q _6885_/A2 _6644_/Z _7750_/Q _7776_/Q _6891_/C1 _6728_/A1 VDD VSS
+ gf180mcu_fd_sc_mcu7t5v0__aoi222_1
X_3936_ _3936_/A1 _3936_/A2 _3936_/A3 _3936_/A4 _3936_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__and4_1
XFILLER_20_810 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_149_366 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3867_ _3886_/A2 hold113/Z _6248_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_4
X_6655_ _7910_/Q _6658_/A2 _6664_/A2 _6891_/B1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor3_4
XFILLER_164_347 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3798_ _7506_/Q _3643_/I hold111/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_5606_ _5735_/A2 _5658_/B _5752_/B1 _5606_/B _5610_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai31_1
X_6586_ _6586_/A1 _6664_/A2 _6586_/B _6587_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_5537_ _5511_/C _5537_/A2 _5739_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_160_520 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_133_712 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_132_211 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_105_425 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5468_ _5031_/B _5473_/A2 _5471_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_87_29 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_7207_ _7961_/Q _7207_/A2 _7207_/B1 _7530_/Q _7207_/C _7208_/A4 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi221_1
X_5399_ _5735_/A2 _5585_/A1 _5724_/B _5759_/A1 _5735_/C _5401_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi221_1
X_4419_ _7979_/Q input88/Z _4420_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__or2_1
X_7138_ _7707_/Q _7190_/C1 _7196_/B1 _7643_/Q _7140_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_7069_ _7778_/Q _7200_/A2 _7200_/B1 _7866_/Q _7075_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_100_152 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_59_567 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_100_174 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2025 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2014 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2003 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_36_33 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2058 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2047 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2036 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1313 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1302 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_54_250 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2069 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1357 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1346 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1335 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1324 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_70_743 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_70_732 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_146_2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1379 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1368 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_167_141 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xinput19 mask_rev_in[23] input19/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_22_191 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_124_701 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_182_177 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_151_520 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_111_428 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_77_73 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_38_707 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_37_228 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_133_90 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_93_50 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_93_83 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_92_389 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_73_570 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_33_434 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_33_445 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1891 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1880 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_4770_ hold680/Z _4773_/A2 _4771_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_174_623 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3721_ _7908_/Q _6585_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__inv_1
XFILLER_173_133 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_173_111 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6440_ hold244/Z _6451_/A2 _6441_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_3652_ _7433_/Q _7001_/C VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_2
XFILLER_173_144 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6371_ _4454_/Z _6383_/A2 _6371_/B _7815_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_61_2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_173_177 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_115_712 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_114_211 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_5322_ _5689_/A2 _5687_/B _5724_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_2
XFILLER_114_233 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_142_575 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5253_ _5689_/A1 _5687_/B _5759_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_4
X_5184_ _5648_/A1 _5752_/B1 _5740_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_4204_ _4204_/A1 _4204_/A2 _4204_/A3 _4204_/A4 _7221_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor4_4
XFILLER_96_673 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4135_ _3835_/Z hold25/Z _5841_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_3_70 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_29_707 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_83_312 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
Xclkbuf_leaf_63_csclk _7961_/CLK _7733_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_56_526 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4066_ _7881_/Q _6503_/A1 _4488_/A1 _7358_/Q _6537_/A1 _7897_/Q _4067_/A4 VDD VSS
+ gf180mcu_fd_sc_mcu7t5v0__aoi222_1
XFILLER_71_507 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_36_250 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_43_209 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_7825_ _7825_/D _7901_/RN _7825_/CLK _7825_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_24_445 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_169_428 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xclkbuf_leaf_78_csclk _7396_/CLK _7510_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_51_264 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_4968_ _5006_/B _5254_/A2 _5709_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_4
X_7756_ _7756_/D _7961_/RN _7756_/CLK _7756_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_51_286 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_52_798 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_4899_ _5006_/B _5006_/C _5392_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_2
XFILLER_149_152 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_137_303 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7687_ _7687_/D _7961_/RN _7735_/CLK _7687_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
X_3919_ _4284_/A1 _7230_/A1 _3921_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_6707_ _6707_/A1 _6767_/C _6707_/B1 _6707_/B2 _7433_/Q _6708_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi221_1
XFILLER_125_7 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_20_673 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6638_ _6878_/A2 _6658_/A2 _6664_/A2 _6893_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor3_4
XFILLER_22_68 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_105_200 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_6569_ _7435_/Q _6622_/A2 _6569_/A3 _6571_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor3_1
XFILLER_145_380 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xclkbuf_leaf_16_csclk _7592_/CLK _7893_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_0_6 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_154_34 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_120_214 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_120_247 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_87_651 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_170_33 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_74_301 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_19_228 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_47_515 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_62_507 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_47_65 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_74_389 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_62_529 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_55_570 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1121 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1132 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1110 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_27_283 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_43_743 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_179_31 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1165 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1154 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1143 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_63_75 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_63_64 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_42_264 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1198 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1187 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1176 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_8_37 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_155_155 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_155_144 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_6_132 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_170_125 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_6_176 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_124_531 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_905 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_916 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_927 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_938 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_949 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_78_673 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_66_802 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_120_770 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5940_ hold633/Z _5953_/A2 _5941_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_18_250 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_179_737 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7610_ _7610_/D _7961_/RN _7694_/CLK _7610_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
X_5871_ _5871_/A1 _7285_/A2 _5873_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_34_776 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_178_247 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4822_ _7498_/Q _4828_/S _4823_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_33_286 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_4753_ hold561/Z _4753_/I1 _4753_/S _7465_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_7541_ _7541_/D _7959_/RN _7545_/CLK hold51/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_147_623 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3704_ _7671_/Q _3704_/ZN VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_7472_ _7472_/D _7961_/RN _7510_/CLK _7472_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
X_4684_ _7465_/Q hold55/Z _4684_/B _4685_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_107_509 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6423_ hold316/Z _6434_/A2 _6424_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_174_486 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_162_648 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_161_114 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3635_ _7554_/Q _3958_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_6354_ _4454_/Z _6366_/A2 _6354_/B _7807_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_108_49 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_5305_ _5682_/A1 _5692_/A2 _5307_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_6285_ hold645/Z _6298_/A2 _6286_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_5236_ _5200_/B _3727_/I _5421_/A1 _5621_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__and3_2
XFILLER_130_534 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_102_225 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_102_236 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_102_214 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_124_37 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5167_ _5735_/A2 _5672_/A2 _5167_/B _5171_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_56_312 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5098_ _5098_/A1 _5098_/A2 _5772_/A1 _5749_/A1 _5106_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand4_1
XFILLER_68_183 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4118_ hold118/Z hold156/Z _4853_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_2
XFILLER_84_676 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4049_ _4049_/A1 _4049_/A2 _4058_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_17_35 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_37_570 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_215 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_204 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_24_242 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_7808_ _7808_/D _7901_/RN _7810_/CLK _7808_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffsnq_1
XPHY_259 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_248 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_237 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_226 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_25_798 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7739_ _7739_/D _7961_/RN _7818_/CLK _7739_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_12_459 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_137_144 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_123_4 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_20_470 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_180_412 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_180_401 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_165_44 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_109_2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_106_531 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_152_169 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_121_567 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xhold8 hold8/I hold8/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
XFILLER_94_429 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_90_602 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_75_698 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_74_41 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_15_231 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_15_286 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_70_392 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_31_757 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_169_792 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_90_84 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_129_689 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
Xhold408 _7682_/Q hold408/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
XFILLER_171_456 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_144_659 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_143_125 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
Xhold419 _7803_/Q hold419/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
XFILLER_7_496 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_152_670 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_112_534 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_97_212 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_97_223 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_713 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_702 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_724 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_6070_ hold68/Z _6072_/A2 _6070_/B hold394/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
XTAP_735 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_746 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_757 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_768 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_39_802 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
Xload_slew344 _7961_/RN _7901_/RN VDD VSS gf180mcu_fd_sc_mcu7t5v0__buf_20
X_5021_ _5529_/A2 _5529_/A3 _5021_/B1 _5010_/Z _5548_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_4
XFILLER_78_481 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_66_621 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_24_2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_779 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_66_676 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_38_378 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_38_389 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_93_495 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6972_ _7798_/Q _7191_/B1 _7201_/B1 _7668_/Q _6972_/C _6976_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi221_1
XFILLER_19_570 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_179_512 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5923_ hold637/Z _5936_/A2 _5924_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_5854_ _7982_/I _5855_/A1 _5855_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_21_212 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_167_718 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4805_ _7224_/I0 _7489_/Q _4809_/S _7489_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_5785_ _5785_/A1 _5795_/A3 _5785_/A3 _5785_/B _5787_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai31_1
X_7524_ _7524_/D _7961_/RN _7650_/CLK _7524_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
X_4736_ hold94/I hold7/Z _4741_/S hold8/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_119_144 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_174_261 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_174_250 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7455_ _7455_/D _7901_/RN _7743_/CLK hold60/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
X_4667_ hold55/Z hold73/Z _4668_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_135_615 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_119_37 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_174_283 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_119_199 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6406_ hold324/Z _6417_/A2 _6407_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_7386_ _7386_/D input75/Z _7391_/CLK _7386_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
X_6337_ _4454_/Z _6349_/A2 _6337_/B _7799_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_4598_ _4454_/Z _4598_/A2 _4598_/B _7402_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_1_628 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_103_567 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6268_ hold663/Z _6281_/A2 _6269_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_5219_ _5452_/C _5543_/C _5545_/A2 _5580_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor3_1
X_6199_ hold415/Z _6208_/A2 _6200_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_76_429 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8007_ _8007_/I _8007_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_151_24 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_151_79 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_57_698 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_60_808 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_44_33 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_157_206 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_52_392 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_12_256 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_9_728 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_126_615 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_165_283 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_109_81 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_109_70 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_79_212 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_39_109 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_48_621 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_85_73 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_48_676 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_75_495 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_90_443 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_63_657 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_50_307 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_50_318 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_176_526 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5570_ _5692_/A1 _5218_/C _5702_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_156_250 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_4521_ hold90/Z _4521_/A2 _4521_/B hold400/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_7240_ _7520_/Q _7240_/A2 _7240_/B1 _7519_/Q _7241_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_4452_ _7506_/Q hold34/Z hold35/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_144_423 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xhold205 _7997_/I hold205/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
Xhold216 hold216/I _7678_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
Xhold249 _7630_/Q hold249/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
Xhold238 hold238/I _6089_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
XFILLER_116_169 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
Xhold227 _7357_/Q hold227/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
XFILLER_171_286 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_131_139 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_113_810 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4383_ _4383_/A1 _4383_/A2 _4383_/B _7413_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_7171_ _7527_/Q _7189_/A2 _7191_/B1 _7405_/Q _7172_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_6122_ hold353/Z _6123_/A2 _6123_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_543 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_532 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_521 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_510 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_6053_ hold68/Z _6055_/A2 _6053_/B hold436/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_86_727 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_85_215 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_554 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_565 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_576 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_5004_ _3722_/I _3723_/I _5254_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_4
XTAP_587 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_598 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_66_473 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_54_602 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_38_175 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_53_112 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_54_646 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1709 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_121_27 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_81_465 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_6955_ _7914_/Q _7913_/Q _6599_/Z _6955_/A4 _7205_/B1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor4_4
X_5906_ hold161/Z hold276/I _5907_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_34_392 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6886_ _6886_/A1 _6886_/A2 _6886_/A3 _6887_/C VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_139_239 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_14_69 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5837_ hold554/Z _5840_/A2 _5838_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_182_507 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5768_ _5122_/Z _5768_/A2 _5768_/A3 _5769_/A4 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_175_570 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_108_615 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_107_103 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4719_ hold108/Z _7285_/A2 _4731_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_4
X_7507_ _7507_/D _7961_/RN _7531_/CLK _7507_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_163_732 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_147_283 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_135_423 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5699_ _5590_/B _5581_/B _5737_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_108_637 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7438_ _7438_/D _7961_/RN _7673_/CLK _7438_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
X_7369_ _7369_/D _7961_/RN _7370_/CLK _7369_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffsnq_2
Xhold761 _7347_/Q hold761/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
XFILLER_1_425 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xhold772 _7644_/Q hold772/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
Xhold750 _7886_/Q hold750/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
XFILLER_150_459 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_150_448 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_162_34 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_130_161 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_89_576 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_77_716 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_39_66 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_130_194 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_176_2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_57_484 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_60_605 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_45_668 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_72_487 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_32_318 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_158_526 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_173_507 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_9_558 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_138_250 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_126_401 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_5_753 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_153_286 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_122_673 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_67_215 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_68_749 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_83_708 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_36_602 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_48_473 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_36_668 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6740_ _7719_/Q _6881_/A2 _6882_/B1 _7655_/Q _6742_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_51_638 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3952_ _7738_/Q _6192_/A1 _6090_/A1 _7690_/Q _3953_/A4 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_16_392 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_91_2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3883_ _3886_/A2 _4075_/B _4232_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_4
X_6671_ _7814_/Q _6880_/A2 _6892_/A2 _7758_/Q _6673_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_5622_ _5622_/A1 _5620_/B _5622_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__or2_1
XFILLER_176_389 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_164_507 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_157_570 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5553_ _5553_/A1 _5553_/A2 _5769_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_145_721 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_129_283 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_8_591 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4504_ hold90/Z _4504_/A2 _4504_/B hold397/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_5484_ _4965_/B _5603_/A1 _5797_/A2 _5485_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor3_1
X_7223_ _7223_/A1 _7228_/S _7223_/B _7944_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_4435_ _7980_/Q input75/Z _4435_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__or2_1
X_4366_ _4366_/A1 _4366_/A2 _4367_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_7154_ _7651_/Q _7195_/A2 _7207_/B1 _7723_/Q _7158_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_6105_ hold343/Z _6106_/A2 _6106_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_113_684 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_98_373 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4297_ _7342_/Q _4308_/S _4296_/Z _4297_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__and3_1
XFILLER_112_194 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_112_183 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_100_312 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_7085_ _7705_/Q _7190_/C1 _7089_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_373 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_384 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_6036_ hold68/Z _6038_/A2 _6036_/B hold383/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
XTAP_395 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_39_440 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2207 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_132_59 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_132_37 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_39_495 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_54_421 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_2229 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2218 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1506 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_82_741 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_13 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
X_7987_ hold97/I _7987_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_1539 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1528 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1517 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_14_318 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_24 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_35 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_46 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_25_35 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_42_605 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_42_638 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_168_802 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6938_ _6938_/I _6948_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XPHY_57 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_68 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_79 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
X_6869_ _7509_/Q _6887_/B1 _6891_/B1 _7507_/Q _6871_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_22_384 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_167_378 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_41_89 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_163_540 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_135_286 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_173_44 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
Xhold580 hold580/I _7471_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
XFILLER_104_673 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xhold591 _7392_/Q hold591/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
XFILLER_103_194 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_49_215 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_49_248 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_65_708 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_18_602 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_18_613 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_122_92 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_122_70 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_60_413 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_17_167 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_32_104 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_45_465 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_159_802 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_60_424 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_32_115 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_33_638 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_139_570 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_127_721 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_181_370 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_154_584 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_142_735 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_141_212 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_141_234 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4220_ _7766_/Q _6265_/A1 _4564_/A1 _7389_/Q _4264_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_4151_ hold275/Z _4151_/A2 _4888_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_110_676 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_95_354 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4082_ _7726_/Q hold119/I _6124_/A1 _7702_/Q _4084_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_68_568 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_95_398 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_7910_ _7910_/D _7961_/RN _7940_/CLK _7910_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffsnq_4
XFILLER_102_18 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7841_ _7841_/D _7901_/RN _7865_/CLK _7841_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_36_443 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_36_454 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_24_605 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4984_ _3723_/I _5777_/A1 _5797_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_2
X_7772_ _7772_/D _7901_/RN _7867_/CLK _7772_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_63_295 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_36_498 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6723_ _7784_/Q _6883_/B1 _6894_/A2 _7840_/Q _6729_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_3935_ input27/Z _4239_/A2 _6537_/A1 _7900_/Q _3936_/A4 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_51_479 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_177_632 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6654_ _6878_/A2 _6658_/A2 _6662_/A3 _6891_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor3_4
XFILLER_177_676 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_176_164 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5605_ _5735_/A2 _5606_/B _5674_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_3866_ hold113/Z hold128/Z _6265_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_4
XFILLER_164_337 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3797_ _7341_/Q _7414_/Q _4303_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_6585_ _7909_/Q _6585_/A2 _6664_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_4
X_5536_ _5543_/B _5153_/C _5536_/A3 _5537_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor3_1
XFILLER_145_562 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_133_702 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5467_ _5602_/A1 _5602_/A2 _5527_/A1 _5473_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor3_1
XFILLER_117_286 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_172_392 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4418_ input83/Z _4418_/I1 _7979_/Q _4418_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_7206_ _7206_/A1 _7206_/A2 _7206_/A3 _7207_/C VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand3_1
X_5398_ _5733_/A2 _5398_/A2 _5586_/A3 _5398_/A4 _5414_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand4_1
XFILLER_160_598 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_113_470 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7137_ _7675_/Q _7201_/B1 _7204_/B1 _7773_/Q _7140_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_98_181 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_86_321 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_59_535 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_4349_ _7902_/Q _6565_/A1 _6622_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_100_142 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_100_120 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7068_ _7068_/A1 _7068_/A2 _7068_/A3 _7068_/A4 _7078_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand4_1
XFILLER_100_164 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6019_ hold68/Z _6021_/A2 _6019_/B hold498/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
XTAP_2015 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2004 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2059 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2048 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2026 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2037 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1314 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1303 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_70_722 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_55_785 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1347 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1336 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1325 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_36_89 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_42_446 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1358 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1369 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_70_788 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_52_33 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_168_33 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_168_676 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_139_2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_128_529 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_10_321 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_182_167 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_182_134 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_170_318 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_151_510 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_123_212 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_2_531 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_151_587 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_151_565 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_117_70 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_96_118 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_2_575 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_2_586 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_93_803 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_77_354 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_93_73 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_45_295 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1870 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_61_766 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_21_619 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1892 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1881 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_3720_ _7909_/Q _6636_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__inv_1
XFILLER_158_164 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_9_141 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_158_175 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3651_ _7905_/Q _6571_/B2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_174_668 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_146_348 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6370_ hold717/Z _6383_/A2 _6371_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_161_318 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5321_ _5724_/B _5648_/B2 _5496_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_54_2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_154_392 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_154_381 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_114_245 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_114_223 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5252_ _5199_/B _5201_/B _3728_/I _5022_/B _5687_/C VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand4_4
XFILLER_115_779 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_142_598 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5183_ _5496_/A1 _5099_/B _5512_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_102_429 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_68_321 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4203_ _4203_/A1 _4203_/A2 _4203_/A3 _4203_/A4 _4204_/A4 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand4_2
X_4134_ hold25/Z _3869_/I _4754_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_68_387 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_56_538 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_113_39 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_83_357 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4065_ _7817_/Q hold134/I _5828_/A1 _7566_/Q _4231_/B1 input67/Z _4067_/A3 VDD VSS
+ gf180mcu_fd_sc_mcu7t5v0__aoi222_1
XFILLER_56_549 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_36_262 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_37_785 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7824_ _7824_/D _7901_/RN _7844_/CLK _7824_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffsnq_1
XFILLER_64_582 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_51_210 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_52_744 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_169_418 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7755_ _7755_/D _7901_/RN _7755_/CLK _7755_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
X_4967_ _3722_/I _3723_/I _5206_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_4
X_4898_ _5006_/B _5006_/C _4898_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__and2_2
X_3918_ _3918_/A1 _3918_/A2 _3917_/Z _7230_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor3_4
X_7686_ _7686_/D _7961_/RN _7694_/CLK _7686_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffsnq_1
X_6706_ _6706_/A1 _6706_/A2 _6706_/A3 _6707_/B2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor3_1
XFILLER_165_624 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_3849_ _3835_/Z hold118/Z _6073_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_4
XFILLER_22_47 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6637_ _7910_/Q _6661_/A3 _6658_/A3 _6880_/C2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor3_4
XFILLER_180_605 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_164_156 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_138_58 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6568_ _7904_/Q _6561_/Z _6570_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_152_318 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_145_370 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5519_ _5519_/A1 _5519_/A2 _5519_/B _5520_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_98_18 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_105_212 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xclkbuf_3_2__f_csclk clkbuf_0_csclk/Z _7396_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
X_6499_ hold427/Z _6502_/A2 _6500_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_154_46 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_105_245 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_87_641 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_86_140 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_75_803 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_59_354 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_59_376 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_47_33 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_90_806 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1122 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1111 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1100 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_27_295 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1155 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1144 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1133 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1199 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1188 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1177 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1166 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_156_602 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_11_641 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_30_449 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_156_646 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_171_627 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_136_370 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_136_392 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_170_159 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_97_416 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_88_62 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_906 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_917 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_111_226 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_111_215 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_97_449 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_928 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_939 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_81_806 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_65_357 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_92_165 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_19_785 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_18_273 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5870_ hold26/Z _4448_/Z hold27/Z hold12/Z _7581_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XFILLER_33_221 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_34_744 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_73_390 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4821_ _7221_/A1 _4828_/S _4821_/B _7497_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
XTAP_2390 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_4752_ hold68/Z _4753_/S _4752_/B _7464_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_7540_ _7540_/D _7959_/RN _7545_/CLK _7540_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_33_298 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_174_410 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4683_ hold55/Z hold90/Z _4684_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_3703_ _7679_/Q _3703_/ZN VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_7471_ _7471_/D _7961_/RN _7531_/CLK _7471_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_162_605 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_119_348 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6422_ _4454_/Z _6434_/A2 _6422_/B _7839_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_3634_ _7555_/Q _4402_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_146_189 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_134_318 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_161_137 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6353_ hold691/Z _6366_/A2 _6354_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_5304_ _5319_/B _5692_/A2 _5307_/B2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_103_716 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6284_ _4448_/Z _6298_/A2 _6284_/B _7774_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_115_598 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_103_738 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5235_ _5685_/B _5292_/B _5614_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_69_641 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_68_140 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5166_ _5643_/A2 _5783_/A2 _5166_/B _5166_/C _5171_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XFILLER_96_460 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_56_302 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_110_270 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_5097_ _5735_/A2 _5669_/A1 _5749_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_4117_ hold113/Z hold107/Z _4574_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_4048_ input55/Z _5886_/A1 _4239_/A2 input23/Z hold26/I _7576_/Q _4049_/A2 VDD VSS
+ gf180mcu_fd_sc_mcu7t5v0__aoi222_1
XFILLER_140_37 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_169_215 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_216 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_205 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_24_254 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_40_703 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_7807_ _7807_/D _7901_/RN _7851_/CLK _7807_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffsnq_1
XPHY_249 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_238 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_227 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
X_5999_ hold514/Z _6004_/A2 _6000_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_178_771 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_138_602 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7738_ _7738_/D _7901_/RN _7818_/CLK _7738_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_33_68 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_40_747 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_177_281 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_149_68 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_20_460 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_149_79 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_138_646 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_138_657 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_138_668 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_137_123 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7669_ _7669_/D _7961_/RN _7701_/CLK _7669_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffsnq_1
XFILLER_180_424 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_153_638 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_118_392 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_79_405 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_161_682 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_133_384 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xoutput290 _7366_/Q pll_trim[3] VDD VSS gf180mcu_fd_sc_mcu7t5v0__buf_8
XFILLER_58_32 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
Xhold9 hold9/I hold9/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
XFILLER_75_655 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_114_93 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_47_357 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_47_379 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_90_636 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_74_176 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_62_316 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_16_744 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_169_771 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_90_41 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_31_747 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_30_268 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_156_443 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_144_605 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xhold409 _7853_/Q hold409/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
XFILLER_116_318 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xclkbuf_leaf_62_csclk clkbuf_opt_1_0_csclk/Z _7692_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_128_189 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_99_50 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_152_693 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_151_170 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_124_362 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_98_747 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xclkbuf_leaf_77_csclk _7396_/CLK _7531_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XTAP_714 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_703 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_725 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_5020_ _5010_/Z _5021_/B1 _5020_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_151_181 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xload_slew345 input75/Z _7961_/RN VDD VSS gf180mcu_fd_sc_mcu7t5v0__buf_20
XTAP_736 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_747 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_758 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_78_460 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_769 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_17_2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_66_666 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_26_508 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6971_ _6971_/A1 _6971_/A2 _6971_/A3 _6972_/C VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_80_135 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_72 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5922_ _4448_/Z _5936_/A2 _5922_/B _7604_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
Xclkbuf_leaf_15_csclk _7592_/CLK _7873_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_110_29 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_80_179 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_61_371 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5853_ hold16/Z hold775/Z hold22/Z _7573_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_5784_ _5784_/A1 _5704_/Z _5784_/A3 _5785_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_61_393 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_22_747 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4804_ _7223_/A1 _4809_/S _4804_/B _7488_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_4735_ hold79/I hold3/Z _4741_/S hold4/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_119_112 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_9_70 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7523_ _7523_/D _7961_/RN _7650_/CLK _7523_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_159_281 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_119_134 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_175_785 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7454_ _7454_/D _7901_/RN _7463_/CLK hold63/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
X_4666_ _7984_/I _4685_/A1 _4669_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_147_465 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_119_167 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_119_156 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_135_638 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6405_ _4454_/Z _6417_/A2 _6405_/B _7831_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_4597_ hold574/Z _4598_/A2 _4598_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_7385_ _7385_/D input75/Z _7391_/CLK _7385_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
X_6336_ hold605/Z _6349_/A2 _6337_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_135_59 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_130_321 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_6267_ _4448_/Z _6281_/A2 _6267_/B _7766_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_139 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5218_ _5421_/B1 _5218_/A2 _5218_/B _5218_/C _5294_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai211_1
X_6198_ _4460_/Z _6208_/A2 _6198_/B hold214/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_8006_ _8006_/I _8006_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_69_460 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_5149_ _5543_/B _5552_/A3 _5548_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_130_398 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_56_121 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_151_58 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_84_463 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_29_357 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_178_6 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_151_69 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_44_327 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_56_176 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_13_769 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_138_443 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_60_33 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_176_33 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_126_605 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_121_2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_176_99 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_153_479 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_125_159 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_134_671 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_121_354 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_48_688 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_141_91 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_90_477 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_62_179 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_62_168 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_172_700 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_157_785 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_156_262 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_117_605 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4520_ hold398/Z _4521_/A2 hold399/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_172_744 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_172_755 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xhold217 _7382_/Q hold217/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
Xhold206 hold206/I _7423_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
XFILLER_117_638 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_116_137 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4451_ hold735/Z _4487_/A1 hold736/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_7_283 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xhold239 hold239/I _7683_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
XFILLER_116_159 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_7_294 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
Xhold228 hold228/I _4494_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
X_7170_ _7521_/Q _7189_/B1 _7189_/C1 _7494_/Q _7172_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_131_107 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_125_682 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_6121_ hold68/Z _6123_/A2 _6121_/B _7698_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_4382_ _4383_/A2 _4382_/A2 _7413_/Q _4383_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
XTAP_500 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_112_321 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_98_566 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_533 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_522 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_511 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_6052_ hold435/Z _6055_/A2 _6053_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_105_29 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_79_780 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_544 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_555 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_566 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_5003_ _5087_/C _5777_/A1 _5741_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_2
XFILLER_112_387 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_577 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_588 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_599 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_39_633 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_66_463 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_26_327 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_53_102 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_81_455 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6954_ _6955_/A4 _6954_/A2 _7205_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_4
X_5905_ _4448_/Z hold276/Z _5905_/B _7596_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_81_499 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_179_354 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_179_343 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6885_ _7505_/Q _6885_/A2 _6885_/B1 _7528_/Q _6886_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_139_229 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_14_37 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_10_717 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_5836_ hold73/Z _5840_/A2 _5836_/B _7566_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_148_741 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5767_ _5331_/Z _5767_/A2 _5767_/A3 _5771_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand3_1
X_7506_ _7506_/D _7959_/RN _7958_/CLK _7506_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_4
XFILLER_147_240 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4718_ _4718_/A1 hold92/Z _4718_/B hold93/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_5698_ _5684_/Z _5698_/A2 _5698_/B _5719_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_108_605 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4649_ hold205/Z _4652_/A1 _4652_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_7437_ _7437_/D _7961_/RN _7689_/CLK _7437_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_116_682 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_104_811 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
Xhold740 _7782_/Q hold740/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
Xhold762 _7355_/Q hold762/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
X_7368_ _7368_/D _7961_/RN _7370_/CLK _7368_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffsnq_1
Xhold751 _7533_/Q hold751/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
Xhold773 _7961_/Q hold773/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
XFILLER_131_641 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6319_ hold729/Z _6332_/A2 _6320_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_1_437 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_7299_ input75/Z _4334_/Z _7299_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_103_376 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_103_354 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_89_588 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_89_599 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_39_45 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_18_806 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_57_463 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_85_783 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_29_165 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_29_176 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_45_636 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_57_496 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_169_2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_72_455 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_72_444 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_17_349 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_44_179 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_111_83 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_111_50 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_71_65 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_13_566 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_139_774 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_154_744 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_154_755 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_126_446 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_113_129 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_5_776 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_106_170 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_96_73 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_492 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_48_463 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_75_282 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_24_809 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3951_ _7714_/Q _6141_/A1 _6158_/A1 _7722_/Q _3953_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_35_157 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_50_105 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_63_499 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_44_680 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3882_ _4075_/B _3881_/Z _4219_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_4
X_6670_ _7644_/Q _6880_/C2 _6644_/Z _7748_/Q _6673_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_5621_ _5624_/A2 _5648_/B2 _5621_/B _5740_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_84_2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5552_ _5543_/B _5153_/C _5552_/A3 _5552_/A4 _5553_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor4_1
XFILLER_129_240 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4503_ hold395/Z _4504_/A2 hold396/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_5483_ _5543_/C _5543_/B _5498_/A2 _5498_/B _5218_/B _5547_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai32_2
XFILLER_6_60 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4434_ _7520_/Q _4338_/Z _7512_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_144_276 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7222_ _7944_/Q _7228_/S _7223_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_4365_ _5224_/A3 _5224_/A4 _4365_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__or2_1
XFILLER_160_747 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_113_641 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_104_129 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7153_ _7153_/A1 _7153_/A2 _7153_/A3 _7153_/A4 _7159_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand4_1
XFILLER_140_460 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7084_ _7753_/Q _7201_/A2 _7201_/B1 _7673_/Q _7100_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_112_151 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6104_ hold68/Z _6106_/A2 _6104_/B _7690_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_86_503 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4296_ _7341_/Q _7340_/Q _4296_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_112_173 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6035_ hold382/Z _6038_/A2 _6036_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_374 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_385 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_396 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2208 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_67_783 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_27_614 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_54_411 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2219 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_7986_ _7986_/I _7986_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
XTAP_1529 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1518 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1507 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_25 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_14 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_36 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_47 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_26_179 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_81_296 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6937_ _6937_/A1 _6954_/A2 _6938_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_4
XPHY_58 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_69 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
X_6868_ _7470_/Q _6659_/Z _6884_/B1 _7521_/Q _6871_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_167_357 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_10_514 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5819_ _4448_/Z _5827_/A2 _5819_/B _7558_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_50_672 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6799_ _6799_/A1 _6799_/A2 _6799_/A3 _6799_/A4 _6799_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__and4_1
XFILLER_182_349 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_108_424 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_151_725 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_173_12 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_1_212 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xhold581 _7508_/Q hold581/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
Xhold570 _7757_/Q hold570/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
Xhold592 _7475_/Q hold592/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
XFILLER_106_50 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_73_720 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_66_76 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_18_625 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_73_764 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_45_444 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_57_282 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_33_628 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_82_53 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_45_499 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_9_312 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_173_327 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_154_530 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_99_105 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_5_562 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_142_747 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_122_460 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_96_812 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4150_ _4153_/A1 _4217_/A2 _4848_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_110_622 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_95_344 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4081_ _7734_/Q _6192_/A1 _6073_/A1 _7678_/Q _6107_/A1 _7694_/Q _4084_/A1 VDD VSS
+ gf180mcu_fd_sc_mcu7t5v0__aoi222_1
XFILLER_49_783 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_7840_ _7840_/D _7901_/RN _7900_/CLK _7840_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffsnq_1
X_4983_ _5206_/A2 _5709_/A1 _5669_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_4
X_7771_ _7771_/D _7901_/RN _7867_/CLK _7771_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_51_425 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6722_ _7377_/Q _6882_/A2 _6712_/Z _6830_/B _6894_/C1 _7832_/Q _6729_/A2 VDD VSS
+ gf180mcu_fd_sc_mcu7t5v0__aoi222_1
X_3934_ _7381_/Q hold114/I _4505_/A1 _7369_/Q _6452_/A1 _7860_/Q _3936_/A3 VDD VSS
+ gf180mcu_fd_sc_mcu7t5v0__aoi222_1
X_3865_ _4212_/A2 hold25/Z _5920_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_4
XFILLER_20_812 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6653_ _6878_/A2 _6663_/A4 _6662_/A3 _6890_/B1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor3_4
XFILLER_149_357 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5604_ _4943_/Z _5604_/A2 _5606_/B _5610_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_176_176 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_117_210 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3796_ hold19/Z _3925_/A2 hold127/Z _3794_/Z _3796_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__or4_4
X_6584_ _6587_/A2 _6584_/A2 _7908_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_5535_ _5535_/A1 _5548_/A3 _5536_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_118_744 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_118_788 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_117_276 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5466_ _5735_/A2 _4996_/Z _5658_/B _5643_/A2 _5674_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_133_769 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_105_449 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_105_438 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7205_ _7534_/Q _7205_/A2 _7205_/B1 _7538_/Q _7206_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_4417_ input84/Z input67/Z _7980_/Q _4417_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_5397_ _5669_/B _5669_/A1 _5292_/B _5621_/B _5583_/B _5398_/A4 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi221_1
XFILLER_87_812 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_141_791 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_7136_ _7781_/Q _7200_/A2 _7203_/B1 _7885_/Q _7140_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_99_694 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_86_300 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4348_ _7902_/Q _6565_/A1 _6622_/A1 _7581_/Q _6572_/A1 _7432_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai32_1
XFILLER_98_193 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_7067_ _7712_/Q _7189_/A2 _7189_/B1 _7688_/Q _7189_/C1 _7656_/Q _7068_/A4 VDD VSS
+ gf180mcu_fd_sc_mcu7t5v0__aoi222_1
XFILLER_47_709 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4279_ _4279_/A1 _4279_/A2 _4279_/A3 _4279_/A4 _4279_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__and4_1
XFILLER_100_176 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_86_388 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6018_ hold497/Z _6021_/A2 _6019_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_27_411 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2016 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2005 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_36_46 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_2049 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2027 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2038 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1304 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_82_550 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_7969_ _7969_/D _7322_/Z _4415_/A2 _7969_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XTAP_1348 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1337 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1326 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1315 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_14_105 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_27_499 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1359 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_11_812 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_128_508 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_10_333 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_22_193 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_168_89 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_167_176 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_136_530 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_10_399 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_6_337 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_136_585 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_124_703 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_124_747 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_108_298 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_123_268 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_96_108 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_104_460 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_131_290 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_77_97 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_38_709 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_18_400 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_133_70 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_58_591 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_61_712 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_93_85 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_33_414 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_33_425 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_159_611 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1860 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_61_778 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_33_447 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1893 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1882 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1871 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_60_266 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_13_160 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_20_108 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_173_113 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3650_ _7904_/Q _6567_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_173_179 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5320_ _5006_/C _5419_/B _5555_/B _5326_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_5251_ _5338_/A1 _5369_/B _5271_/A3 _5624_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor3_4
XFILLER_142_522 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_114_268 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_69_812 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_47_2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4202_ _4202_/A1 _4202_/A2 _4202_/A3 _4203_/A4 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor3_1
XFILLER_123_780 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5182_ _5797_/B _5797_/C _5741_/A3 _5185_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor3_1
XFILLER_95_130 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_95_141 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_84_804 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_29_709 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4133_ hold118/Z _4155_/A2 _4858_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_2
XFILLER_110_463 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4064_ _7607_/Q _5920_/A1 _4505_/A1 _7366_/Q _6005_/A1 _7647_/Q _4067_/A2 VDD VSS
+ gf180mcu_fd_sc_mcu7t5v0__aoi222_1
XFILLER_28_208 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_113_29 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_36_274 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_52_734 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_7823_ _7823_/D _7901_/RN _7895_/CLK _7823_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffsnq_1
X_7754_ _7754_/D _7901_/RN _7755_/CLK _7754_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_24_447 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_149_110 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_4966_ _5309_/A1 _5087_/C _4969_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_6705_ _6705_/A1 _6705_/A2 _6705_/A3 _6705_/A4 _6706_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand4_1
XFILLER_177_441 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3917_ _3917_/A1 _3917_/A2 _3917_/A3 _3917_/A4 _3917_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__or4_1
X_7685_ _7685_/D _7961_/RN _7815_/CLK _7685_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffsnq_1
X_4897_ _4454_/Z _4897_/A2 _4897_/B _7538_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_177_496 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_165_614 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_165_636 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3848_ hold118/Z hold128/Z _6141_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_4
XFILLER_22_37 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_6636_ _6636_/A1 _7908_/Q _6658_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_4
XFILLER_138_37 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_118_530 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3779_ _7977_/Q hold11/I _3780_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_6567_ _6567_/A1 _6565_/B _6567_/B1 _6557_/I _7904_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai22_1
XFILLER_164_179 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5518_ _5547_/A1 _5518_/A2 _5518_/A3 _5519_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor3_1
XFILLER_106_747 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6498_ hold47/Z _6502_/A2 _6498_/B _7875_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_5449_ _5714_/A1 _5797_/A2 _5543_/C _5452_/C _5450_/C VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XFILLER_78_108 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_7119_ _7650_/Q _7195_/A2 _7195_/B1 _7626_/Q _7195_/C1 _7876_/Q _7121_/A3 VDD VSS
+ gf180mcu_fd_sc_mcu7t5v0__aoi222_1
XFILLER_74_303 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_101_496 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_74_325 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_62_509 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_55_561 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_103_73 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_1123 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1112 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1101 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_63_33 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_15_425 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_15_436 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_28_797 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_42_211 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_43_712 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_43_745 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xclkbuf_1_1__f_wbbd_sck clkbuf_0_wbbd_sck/Z _3666__1/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_151_2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1156 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_70_553 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_1145 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1134 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1189 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1178 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1167 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_168_463 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_10_185 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_170_105 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_155_168 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_109_585 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_109_596 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_163_190 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_2_340 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_907 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_112_739 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_97_428 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_918 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_929 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_120_761 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_77_141 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_19_764 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_92_199 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_33_211 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2380 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_179_739 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4820_ _7497_/Q _4828_/S _4821_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_2391 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_21_428 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_33_277 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4751_ hold255/Z _4753_/S _4752_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_1
XTAP_1690 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_159_496 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_147_636 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4682_ hold97/Z _4685_/A1 hold98/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_3702_ _7687_/Q _3702_/ZN VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_7470_ _7470_/D _7961_/RN _7627_/CLK _7470_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
X_3633_ _7973_/Q _3765_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_6421_ hold688/Z _6434_/A2 _6422_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_146_179 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6352_ _4448_/Z _6366_/A2 _6352_/B _7806_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_108_29 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5303_ _3728_/I _5022_/B _5303_/A3 _5303_/A4 _5692_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand4_4
XFILLER_142_341 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_115_566 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6283_ hold739/Z _6298_/A2 _6284_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_142_385 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5234_ _5687_/B _5365_/B1 _5292_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_4
XFILLER_102_205 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5165_ _5006_/B _5206_/A2 _5476_/B _5319_/C _5692_/B _5645_/A1 _5166_/C VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai33_1
XFILLER_111_783 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_110_260 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_69_697 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4116_ hold113/Z hold156/Z _4522_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_96_483 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_96_494 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5096_ _5669_/A1 _5783_/A2 _5772_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_83_122 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_4047_ _7378_/Q hold114/I _4444_/A1 _7350_/Q _6333_/A1 _7801_/Q _4049_/A1 VDD VSS
+ gf180mcu_fd_sc_mcu7t5v0__aoi222_1
XFILLER_83_144 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_71_339 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_25_712 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7806_ _7806_/D _7901_/RN _7806_/CLK _7806_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffsnq_1
XPHY_206 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_52_531 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_52_553 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_239 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_228 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_217 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
X_5998_ hold41/Z _6004_/A2 _5998_/B hold367/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_52_564 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_4949_ _4951_/B _4979_/A3 _5458_/C VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_2
X_7737_ _7737_/D _7901_/RN _7818_/CLK _7737_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_137_102 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7668_ _7668_/D _7961_/RN _7733_/CLK _7668_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffsnq_1
X_6619_ _7918_/Q _6621_/A2 _6620_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_153_628 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_152_105 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7599_ _7599_/D _7901_/RN _7673_/CLK _7599_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_4_605 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_165_499 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_165_46 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_180_469 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_133_352 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_106_566 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_3_148 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_79_428 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
Xoutput280 _7349_/Q pll_trim[18] VDD VSS gf180mcu_fd_sc_mcu7t5v0__buf_8
XFILLER_0_811 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_121_558 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_121_547 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
Xoutput291 _7367_/Q pll_trim[4] VDD VSS gf180mcu_fd_sc_mcu7t5v0__buf_8
XFILLER_58_99 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_74_122 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_114_83 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_74_166 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_74_43 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_62_328 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_130_82 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_43_597 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_169_783 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_156_400 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_129_636 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_30_247 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_30_258 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_156_455 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_128_179 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_7_454 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_171_425 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_99_73 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_140_812 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_124_374 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_3_682 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_715 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_704 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_124_396 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_726 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_737 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_748 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_759 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_120_591 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_120_580 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_78_494 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_93_442 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6970_ _7862_/Q _7200_/B1 _7205_/B1 _7740_/Q _6971_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_65_144 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_65_177 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5921_ hold747/Z _5936_/A2 _5922_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_34_531 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5852_ hold21/Z _7285_/A2 hold22/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_167_709 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5783_ _5104_/B _5783_/A2 _5783_/B _5783_/C _5784_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi211_1
X_4803_ _7488_/Q _4809_/S _4804_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_4734_ _7450_/Q hold16/Z _4741_/S hold17/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_7522_ _7522_/D _7961_/RN _7532_/CLK _7522_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_119_124 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4665_ _4685_/A1 _4665_/A2 _4665_/B hold56/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_134_105 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7453_ _7453_/D _7901_/RN _7461_/CLK hold82/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_147_499 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_134_116 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_7384_ _7384_/D _7901_/RN _7398_/CLK _7384_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
X_4596_ _4448_/Z _4598_/A2 _4596_/B _7401_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_6404_ hold657/Z _6417_/A2 _6405_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_143_661 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6335_ _4448_/Z _6349_/A2 _6335_/B _7798_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_142_171 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_131_812 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_103_503 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_107 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_88_247 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_8005_ _8005_/I _8005_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_6266_ hold730/Z _6281_/A2 _6267_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_5217_ _5392_/A1 _5254_/A3 _5218_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_130_377 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_6197_ hold212/Z _6208_/A2 hold213/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_69_472 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5148_ _5369_/B _5040_/B _5552_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_97_792 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_69_483 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_29_314 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5079_ _5087_/B _5456_/A2 _5079_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_57_678 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_71_114 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_12_203 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_25_586 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_44_57 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_13_759 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_9_708 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_40_534 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_12_247 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_100_74 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_181_712 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_176_56 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_138_455 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_126_617 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_153_425 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_114_2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_109_83 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_106_341 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_140_108 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_122_812 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_95_707 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_663 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_674 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_85_31 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_47_144 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_63_637 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_62_103 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_35_306 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_141_70 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_16_531 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_43_361 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_149_709 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_31_534 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_31_545 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_31_556 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_31_567 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_157_753 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_129_422 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_8_741 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_8_763 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_129_499 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_116_105 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xhold207 _7670_/Q hold207/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
X_4450_ _4487_/A1 _4448_/Z _4450_/B _7347_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
Xhold218 _7667_/Q hold218/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
Xhold229 hold229/I _7357_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
X_4381_ _7965_/Q _7964_/Q _4327_/S _3738_/Z _4383_/A1 _7414_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai32_1
XFILLER_113_812 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6120_ hold401/Z _6123_/A2 _6121_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_98_534 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_534 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_523 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_512 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_501 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_6051_ hold47/Z _6055_/A2 _6051_/B hold296/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
XTAP_545 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_556 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_567 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_5002_ _3723_/I _5662_/A1 _5643_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_4
XFILLER_85_228 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_578 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_589 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_93_272 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_81_423 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_38_188 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_39_689 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_26_339 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6953_ _6953_/A1 _6953_/A2 _6955_/A4 _7202_/B1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor3_4
X_5904_ hold164/Z hold276/I _5905_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_6884_ _7372_/Q _6644_/Z _6884_/B1 _7522_/Q _6886_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_5835_ hold488/Z _5840_/A2 _5836_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_22_534 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5766_ _5766_/A1 _5766_/A2 _5766_/A3 _5767_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor3_1
XFILLER_163_712 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_148_764 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_147_230 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4717_ _7603_/Q _3819_/Z hold91/Z hold92/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_5697_ _5419_/B _5697_/A2 _5697_/A3 _5697_/A4 _5698_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor4_1
X_7505_ _7505_/D _7961_/RN _7871_/CLK _7505_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_162_211 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4648_ _4652_/A1 _4648_/A2 _4648_/B hold198/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_135_425 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_107_116 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_7436_ _7436_/D _7961_/RN _7689_/CLK _7436_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_30_37 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_146_37 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xhold730 _7766_/Q hold730/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
XFILLER_122_108 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
Xhold741 _7798_/Q hold741/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
Xhold763 _7363_/Q hold763/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
X_7367_ _7367_/D _7961_/RN _7587_/CLK _7367_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffsnq_2
Xhold752 _7523_/Q hold752/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
X_4579_ _4579_/A1 _7285_/A2 _4583_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_7298_ _7901_/RN _4334_/Z _7298_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_131_631 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6318_ _4448_/Z _6332_/A2 _6318_/B _7790_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
Xhold774 _7558_/Q hold774/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
XFILLER_130_152 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_130_141 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_89_567 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6249_ hold748/Z _6264_/A2 _6250_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_29_144 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_57_442 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_84_250 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xclkbuf_leaf_61_csclk clkbuf_opt_2_0_csclk/Z _7706_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_29_155 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_111_73 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_111_95 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_71_33 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_9_516 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_9_505 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
Xclkbuf_leaf_76_csclk _7396_/CLK _7627_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_13_578 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_40_386 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_166_550 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_166_594 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_181_531 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_141_428 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_107_661 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_153_299 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_134_480 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xclkbuf_leaf_14_csclk _7592_/CLK _7883_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_136_81 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_122_664 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_121_141 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_67_239 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
Xhold90 hold90/I hold90/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
XFILLER_152_80 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
Xclkbuf_leaf_29_csclk _7825_/CLK _7805_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_75_250 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_90_220 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3950_ _7626_/Q _5954_/A1 _6073_/A1 _7682_/Q _4176_/C _3953_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi221_2
XFILLER_177_804 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3881_ hold19/Z _3925_/A2 hold127/Z _3963_/A4 _3881_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__or4_2
XFILLER_31_353 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5620_ _5681_/A1 _5722_/A1 _5620_/B _5632_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_5551_ _5644_/A2 _5739_/A2 _5551_/A3 _5557_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_77_2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_172_520 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_145_712 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_144_211 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_144_200 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_8_582 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4502_ hold68/Z _4504_/A2 _4502_/B hold537/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_172_531 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5482_ _5648_/A1 _5608_/B _5648_/B2 _5482_/B2 _5644_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_117_469 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7221_ _7221_/A1 _7228_/S _7221_/B _7943_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_172_575 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_104_119 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_104_108 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4433_ _7587_/Q input39/Z _4433_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__and2_1
X_4364_ _5224_/A3 _5224_/A4 _5302_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_2
X_7152_ _7797_/Q _7190_/A2 _7196_/A2 _7893_/Q _7153_/A4 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_4295_ _7339_/Q _4294_/Z _4308_/S VDD VSS gf180mcu_fd_sc_mcu7t5v0__and2_1
X_6103_ hold377/Z _6106_/A2 _6104_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_7083_ _7936_/Q _7133_/S _7109_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_6034_ hold47/Z _6038_/A2 _6034_/B hold405/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
XTAP_375 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_112_196 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_86_559 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_397 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_386 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_66_250 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2209 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_7985_ _7985_/I _7985_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_82_732 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1519 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1508 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_6936_ _6936_/A1 _6936_/A2 _6954_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_2
XPHY_26 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_15 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_37 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_81_286 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_48 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_25_37 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_59 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_41_128 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_179_141 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6867_ _6867_/A1 _6867_/A2 _6867_/A3 _6867_/A4 _6867_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__and4_1
X_6798_ _7843_/Q _6894_/A2 _6659_/Z _7625_/Q _6890_/B1 _7851_/Q _6799_/A4 VDD VSS
+ gf180mcu_fd_sc_mcu7t5v0__aoi222_1
XFILLER_10_504 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5818_ hold774/Z _5827_/A2 _5819_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_50_695 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5749_ _5749_/A1 _5749_/A2 _5749_/A3 _5749_/A4 _5754_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand4_1
XFILLER_182_317 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_41_69 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_136_767 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_136_756 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_135_222 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_123_428 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7419_ hold84/Z _7901_/RN _7461_/CLK _7993_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
Xhold560 _4741_/Z _7457_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
XFILLER_150_247 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_104_620 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_2_747 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xhold571 _7390_/Q hold571/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
XFILLER_103_141 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_1_235 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
Xhold593 hold593/I _7475_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
Xhold582 hold582/I _4847_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
XFILLER_104_697 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_103_185 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_103_152 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_77_515 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_66_44 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_66_33 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_181_2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_85_570 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_64_209 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_82_32 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_72_242 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_17_169 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_72_275 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_14_810 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_15_70 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_9_357 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_127_712 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_154_542 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_181_372 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_147_80 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_181_383 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_141_269 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_68_504 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_122_472 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_110_601 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_68_548 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_68_526 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_1_780 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4080_ _4080_/A1 _4080_/A2 _4080_/A3 _4107_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand3_2
XFILLER_48_250 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_63_264 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4982_ _3722_/I _5006_/B _5254_/A2 _5662_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand3_4
X_7770_ _7770_/D _7901_/RN _7897_/CLK _7770_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_64_798 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_63_286 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_23_106 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_51_415 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3933_ _7876_/Q _6486_/A1 _6022_/A1 _7658_/Q _3936_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_6721_ _7694_/Q _6881_/B1 _6721_/B _6721_/C _6729_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XFILLER_32_651 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_51_459 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3864_ _3801_/Z _3864_/A2 hold24/Z hold274/I hold25/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand4_4
X_6652_ _7838_/Q _6894_/A2 _6887_/B1 _7676_/Q _6683_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_32_673 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5603_ _5603_/A1 _4993_/B _5753_/A2 _5798_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor3_1
XFILLER_31_172 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_176_188 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3795_ _3801_/S hold154/Z _3795_/B _3963_/A4 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi21_4
XFILLER_118_734 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6583_ _7908_/Q _6586_/A1 _6586_/B _6584_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand3_1
X_5534_ _5752_/C _5534_/A2 _5534_/A3 _5644_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor3_1
X_5465_ _5465_/A1 _5803_/A1 _5772_/A3 _5799_/A1 _5472_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand4_1
X_4416_ _3810_/S _4416_/A2 _5903_/A2 _4416_/B2 _4416_/ZN VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai22_1
XFILLER_160_534 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_132_236 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_105_428 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7204_ _7400_/Q _7204_/A2 _7204_/B1 _7390_/Q _7208_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_132_247 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5396_ _5585_/A1 _5672_/A2 _5624_/B _5759_/A1 _5586_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_7135_ _7001_/C _7937_/Q _7161_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_4347_ _7903_/Q _4347_/A2 _4360_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_100_133 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_86_356 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4278_ _7878_/Q _6503_/A1 hold108/I input61/Z _4279_/A4 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_7066_ _7898_/Q _7197_/A2 _7196_/A2 _7890_/Q _7196_/B1 _7640_/Q _7068_/A3 VDD VSS
+ gf180mcu_fd_sc_mcu7t5v0__aoi222_1
XFILLER_74_518 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_67_570 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6017_ hold47/Z _6021_/A2 _6017_/B hold513/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
XTAP_2006 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_39_283 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2039 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2017 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2028 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1305 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_54_242 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_7968_ _7968_/D _7321_/Z _4415_/A2 _7968_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
Xclkbuf_1_0__f_wbbd_sck clkbuf_0_wbbd_sck/Z net299_2/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XTAP_1338 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1327 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1316 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_54_264 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_54_275 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7899_ _7899_/D _7901_/RN _7899_/CLK _7899_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XTAP_1349 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_6919_ _7914_/Q _7913_/Q _6950_/A1 _6941_/A2 _7195_/B1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor4_4
XFILLER_52_46 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_167_144 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_23_695 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_109_712 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_108_211 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_10_389 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_136_575 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_124_759 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_151_567 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_117_61 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_117_50 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_104_450 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xhold390 _7448_/Q hold390/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
XFILLER_7_2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_151_589 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_89_150 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_77_32 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_2_577 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_93_805 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_73_562 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_93_97 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_45_286 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_46_798 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1861 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1850 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_159_634 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1894 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1883 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1872 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_14_673 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_173_103 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_142_534 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5250_ _5779_/A1 _5425_/B _5783_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_114_225 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_114_247 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4201_ _4201_/A1 _4201_/A2 _4202_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_5181_ _5648_/A1 _5066_/Z _5608_/B _5186_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_96_610 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_68_323 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_68_345 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4132_ _4075_/B hold128/Z _5812_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_3_73 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_96_676 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4063_ _4063_/A1 _4063_/A2 _4063_/A3 _4063_/A4 _4068_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand4_1
XFILLER_68_389 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_49_570 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_56_518 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_37_776 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_7822_ _7822_/D _7901_/RN _7834_/CLK _7822_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffsnq_1
XFILLER_51_212 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7753_ _7753_/D _7901_/RN _7753_/CLK _7753_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
X_4965_ _5797_/B _5363_/A2 _4965_/B _4969_/C VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi21_2
XFILLER_51_223 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3916_ _3916_/A1 _3916_/A2 _3916_/A3 _3916_/A4 _3917_/A4 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand4_1
X_6704_ _7749_/Q _6644_/Z _6884_/B1 _7685_/Q _6705_/A4 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_149_144 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7684_ _7684_/D _7961_/RN _7692_/CLK _7684_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffsnq_1
X_4896_ hold686/Z _4897_/A2 _4897_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_3847_ hold123/Z _3787_/Z hold127/Z _3794_/Z _3847_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__or4_4
XFILLER_20_676 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_22_27 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_6635_ _6878_/A2 _6664_/A2 _6661_/A3 _6883_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor3_4
XFILLER_138_49 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6566_ _6567_/A1 _6561_/Z _6567_/B1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_3778_ _3778_/I _7964_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_145_361 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5517_ _5517_/A1 _5642_/A3 _5517_/A3 _5517_/A4 _5518_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand4_1
XFILLER_4_809 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6497_ hold448/Z _6502_/A2 _6498_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_154_37 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5448_ _5448_/A1 _5777_/A2 _5448_/B _5461_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_133_567 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5379_ _5714_/A1 _5689_/A1 _5543_/C _5452_/C _5380_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi211_2
X_7118_ _7698_/Q _7194_/A2 _7194_/B1 _7666_/Q _7194_/C1 _7812_/Q _7121_/A2 VDD VSS
+ gf180mcu_fd_sc_mcu7t5v0__aoi222_1
XFILLER_101_442 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_75_805 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_59_334 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_59_323 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_7049_ _7777_/Q _7200_/A2 _7193_/B1 _7631_/Q _7053_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_47_35 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_47_507 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_86_197 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_28_743 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_70_510 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1113 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1102 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_27_286 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_82_392 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1146 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1124 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1135 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_144_2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1179 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1168 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1157 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_11_698 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_7_636 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_6_124 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_164_681 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_124_534 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_124_523 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_124_512 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_6_179 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_2_330 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_908 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_919 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_93_602 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_78_676 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_65_304 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_80_318 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_61_521 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_61_510 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2370 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2392 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2381 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_4750_ hold627/Z _4750_/I1 _4753_/S _7463_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XTAP_1691 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1680 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_4681_ _4685_/A1 hold69/Z _4681_/B hold70/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_119_328 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_3701_ _7695_/Q _3701_/ZN VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_146_147 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3632_ _7975_/Q _3760_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_6420_ _4448_/Z _6434_/A2 _6420_/B _7838_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_6351_ hold642/Z _6366_/A2 _6352_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_5302_ _5302_/A1 _5011_/B _5302_/A3 _5319_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand3_4
XFILLER_155_692 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_115_534 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_115_545 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6282_ _6282_/A1 _7285_/A2 _6298_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_4
XFILLER_170_695 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_170_673 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5233_ _5254_/A2 _5616_/A1 _5365_/B1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_2
XFILLER_103_718 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5164_ _4993_/C _5452_/C _5543_/C _5559_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor3_1
XFILLER_124_29 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_68_131 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_111_773 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_110_250 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_84_602 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4115_ hold133/Z _4155_/A2 _7285_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_57_805 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5095_ _5669_/A1 _5658_/B _5608_/B _4996_/Z _5095_/C _5098_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi221_1
X_4046_ _4046_/A1 _4046_/A2 _4046_/A3 _4046_/A4 _4058_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand4_1
XFILLER_140_28 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_7805_ _7805_/D _7901_/RN _7805_/CLK _7805_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XPHY_207 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_64_392 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_229 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_218 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
X_5997_ hold366/Z _6004_/A2 _5998_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_4948_ _4944_/Z _4955_/A2 _5741_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_4
X_7736_ _7736_/D _7901_/RN _7819_/CLK _7736_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
X_7667_ _7667_/D _7901_/RN _7806_/CLK _7667_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
X_4879_ hold681/Z _4882_/A2 _4880_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_177_283 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_138_648 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6618_ _7435_/Q _7433_/Q _6618_/A3 _6618_/B _6621_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai31_1
XFILLER_165_478 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_116_6 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7598_ _7598_/D _7901_/RN _7691_/CLK _7598_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_146_692 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_106_534 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6549_ hold47/Z _6553_/A2 _6549_/B _7899_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_118_394 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_161_684 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_160_172 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_160_150 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
Xoutput270 _7565_/Q pll_sel[2] VDD VSS gf180mcu_fd_sc_mcu7t5v0__buf_8
Xoutput281 _7350_/Q pll_trim[19] VDD VSS gf180mcu_fd_sc_mcu7t5v0__buf_8
Xoutput292 _7368_/Q pll_trim[5] VDD VSS gf180mcu_fd_sc_mcu7t5v0__buf_8
XFILLER_58_34 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_75_602 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_59_153 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_48_805 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_58_89 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_114_51 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_101_283 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_87_495 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_74_112 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_101_294 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_90_605 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_75_657 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_74_33 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_90_616 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_90_627 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_90_638 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_62_318 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_15_212 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_28_595 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_43_532 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_90_43 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_168_250 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_128_103 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_128_114 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_23_70 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_156_467 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_7_444 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_143_139 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_125_810 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_7_499 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_99_85 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_152_662 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_97_215 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_716 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_705 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_727 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_738 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_749 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_66_602 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_93_410 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_78_473 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_171_90 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_93_454 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_19_551 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_41 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5920_ _5920_/A1 hold32/Z _5936_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_4
XFILLER_46_392 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_179_548 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_22_727 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5851_ _4448_/Z _5851_/A2 _5851_/B _7572_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_179_559 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5782_ _5782_/A1 _5782_/A2 _5782_/A3 _5795_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_21_215 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4802_ _7221_/A1 _4809_/S _4802_/B _7487_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_4733_ _3830_/Z _4742_/A2 _4741_/S VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_4
X_7521_ _7521_/D _7961_/RN _7642_/CLK _7521_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_159_283 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7452_ hold8/Z _7901_/RN _7461_/CLK hold94/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_9_94 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4664_ hold9/Z hold55/Z _4664_/B _4665_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_119_29 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6403_ _4448_/Z _6417_/A2 _6403_/B _7830_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_7383_ _7383_/D _7901_/RN _7802_/CLK _7383_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
X_4595_ hold656/Z _4598_/A2 _4596_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_89_705 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6334_ hold741/Z _6349_/A2 _6335_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_6265_ _6265_/A1 _7285_/A2 _6281_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_4
XFILLER_88_204 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5216_ _5200_/B _3727_/I _5369_/B _5421_/B1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand3_2
X_8004_ _8004_/I _8004_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_6196_ _4454_/Z _6208_/A2 _6196_/B _7733_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_5147_ _5528_/A2 _5020_/Z _5153_/C VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_2
XFILLER_130_389 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_111_570 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_69_495 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_28_37 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_29_304 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_57_635 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5078_ _3722_/I _5392_/A1 _5456_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_2
XFILLER_72_605 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_178_8 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4029_ input48/Z _4275_/A2 _5920_/A1 _7608_/Q _4030_/A4 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_44_318 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_71_126 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_13_716 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_25_576 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_25_565 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_52_362 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_40_513 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_52_373 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7719_ _7719_/D _7901_/RN _7821_/CLK _7719_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_21_771 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_166_798 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_165_286 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_109_73 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_107_2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_161_470 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_134_673 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_133_150 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_109_95 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_79_215 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_87_281 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_47_134 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_85_87 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_35_318 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_62_126 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_28_392 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_71_671 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_43_340 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_70_170 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_169_570 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_129_434 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_12_771 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_129_478 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_79_6 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_7_230 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_171_212 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xhold208 hold208/I _7670_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
Xhold219 hold219/I _6055_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
XFILLER_116_139 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_109_191 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4380_ _4292_/B _4380_/A2 _4380_/B _7415_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_113_802 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_112_312 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_524 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_513 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_502 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_6050_ hold295/Z _6055_/A2 _6051_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_140_676 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_112_345 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_79_771 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_546 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_535 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_557 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_112_389 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5001_ _5600_/A1 _5363_/A2 _5663_/A1 _5585_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor3_2
XTAP_568 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_579 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_22_2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_66_454 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_94_796 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_26_318 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_38_167 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_54_605 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_121_19 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_93_295 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_6952_ _6953_/A1 _6599_/Z _6955_/A4 _7204_/B1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor3_4
XFILLER_179_323 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5903_ _5903_/A1 _5903_/A2 hold32/Z hold276/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand3_4
X_6883_ _7406_/Q _6883_/A2 _6883_/B1 _7398_/Q _6886_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_179_345 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_61_170 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5834_ _4460_/Z _5840_/A2 _5834_/B hold157/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_22_524 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_167_507 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5765_ _5765_/A1 _5765_/A2 _5765_/A3 _5766_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand3_1
X_4716_ _3819_/Z hold90/Z hold91/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_5696_ _5686_/Z _5696_/A2 _5695_/Z _5697_/A4 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand3_1
X_7504_ _7504_/D _7961_/RN _7587_/CLK _7504_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
X_4647_ _7456_/Q _3830_/Z _4647_/B _4648_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_147_286 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_135_437 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7435_ _7435_/D _7961_/RN _7940_/CLK _7435_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_2
X_7366_ _7366_/D _7961_/RN _7565_/CLK _7366_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffsnq_2
Xhold720 _7391_/Q hold720/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
XFILLER_162_267 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
Xhold753 _7341_/Q hold753/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
XFILLER_116_673 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_100_9 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_89_513 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
Xhold731 _7854_/Q hold731/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
X_6317_ hold745/Z _6332_/A2 _6318_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
Xhold742 _7822_/Q hold742/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
Xhold764 _7569_/Q hold764/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
X_4578_ _4454_/Z _4578_/A2 _4578_/B _7394_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_7297_ _7901_/RN _4334_/Z _7297_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_143_492 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_103_312 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_89_535 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_1_428 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xhold775 _7573_/Q hold775/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
X_6248_ _6248_/A1 hold32/Z _6264_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_4
X_6179_ _4454_/Z _6191_/A2 _6179_/B _7725_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_162_37 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_29_101 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_69_281 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_57_432 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_85_785 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_85_774 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_72_402 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_29_167 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_44_104 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_45_605 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_45_638 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_72_479 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_111_41 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_25_373 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_52_170 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_71_23 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_40_321 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_40_376 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_40_398 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_153_212 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_5_712 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_181_576 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_113_109 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_107_651 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_4_266 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_122_676 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_121_120 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_96_75 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_95_516 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_96_97 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
Xhold80 hold80/I hold80/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
Xhold91 hold91/I hold91/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
XFILLER_36_605 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_91_755 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_75_295 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_63_446 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_63_424 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_90_243 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_44_660 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3880_ hold275/Z _3835_/Z _6469_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_4
XFILLER_43_192 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_176_337 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_5550_ _5179_/B _5672_/A2 _5550_/B _5550_/C _5551_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XFILLER_172_510 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_129_286 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_129_275 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5481_ _5658_/B _5179_/B _5757_/B _5765_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_4501_ hold535/Z _4504_/A2 hold536/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_7220_ _7943_/Q _7228_/S _7221_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_4432_ _7586_/Q input70/Z _4432_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__and2_1
X_4363_ _5302_/A1 _5195_/B _4906_/S VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_2
XFILLER_153_790 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_125_492 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_125_470 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7151_ _7691_/Q _7189_/B1 _7189_/C1 _7659_/Q _7153_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_98_321 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4294_ _7338_/Q _7337_/Q _7336_/Q _4294_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__and3_1
XFILLER_113_643 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6102_ hold47/Z _6106_/A2 _6102_/B _7689_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_86_505 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7082_ _7133_/S _7082_/A2 _7082_/B _7935_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_6033_ hold404/Z _6038_/A2 _6034_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_58_207 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_376 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_100_337 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_398 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_387 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_132_29 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_66_240 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_7984_ _7984_/I _7984_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_27_638 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1509 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_82_788 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_81_243 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_27 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_16 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_38 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_25_27 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_6935_ _6941_/A2 _6935_/A2 _7190_/C1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_4
XPHY_49 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_22_321 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6866_ _7371_/Q _6644_/Z _6665_/Z _7537_/Q _6891_/C1 _7393_/Q _6867_/A4 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi222_1
XFILLER_167_348 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6797_ _7795_/Q _6893_/A2 _6893_/B1 _7771_/Q _6893_/C1 _7633_/Q _6799_/A3 VDD VSS
+ gf180mcu_fd_sc_mcu7t5v0__aoi222_1
X_5817_ _5817_/A1 _7285_/A2 _5827_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_4
XFILLER_148_551 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5748_ _5748_/A1 _5748_/A2 _5777_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__or2_1
X_5679_ _5679_/A1 _5679_/A2 _5698_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_7418_ hold96/Z _7901_/RN _7461_/CLK _7992_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
Xhold561 _7465_/Q hold561/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
XFILLER_9_6 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
Xhold550 hold550/I _7366_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
Xhold572 _7534_/Q hold572/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
X_7349_ _7349_/D _7961_/RN _7570_/CLK _7349_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffsnq_2
XFILLER_103_120 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_89_354 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xhold583 hold583/I _7508_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
Xhold594 _7887_/Q hold594/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
XFILLER_104_676 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_77_527 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_58_752 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_18_605 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_174_2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_85_593 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_85_582 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_72_232 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_45_479 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_26_693 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_41_641 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_13_354 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_139_540 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_41_696 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_127_702 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_166_392 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_31_70 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_147_70 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_126_256 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_141_226 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_141_215 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_122_451 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_68_538 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_95_357 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_95_335 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_64_744 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_63_221 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_36_435 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_48_295 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_91_563 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_91_552 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4981_ _5309_/A1 _5709_/A1 _5777_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_4
XFILLER_91_585 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_3932_ _7730_/Q hold119/I _6124_/A1 _7706_/Q _6107_/A1 _7698_/Q _3936_/A1 VDD VSS
+ gf180mcu_fd_sc_mcu7t5v0__aoi222_1
X_6720_ _6720_/A1 _6720_/A2 _6720_/A3 _6721_/C VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_177_624 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_3863_ _4075_/B _4151_/A2 _4249_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_4
XFILLER_31_140 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6651_ _7910_/Q _6664_/A2 _6661_/A3 _6887_/B1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor3_4
X_5602_ _5602_/A1 _5602_/A2 _5797_/A2 _5602_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__or3_1
X_6582_ _7434_/Q _6585_/A2 _6590_/A1 _6587_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_164_329 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_164_318 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5533_ _5533_/A1 _5543_/B _5153_/C _5552_/A4 _5534_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor4_1
X_3794_ hold104/Z hold154/Z _3801_/S _3794_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_4
XFILLER_145_521 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_117_223 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_117_212 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_11_29 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_127_29 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5464_ _5669_/B _5643_/A2 _5608_/B _4996_/Z _5799_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_1
Xclkbuf_leaf_60_csclk clkbuf_3_6__f_csclk/Z _7702_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
X_4415_ _3810_/S _4415_/A2 _4416_/B2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_132_215 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5395_ _5669_/A1 _5783_/A2 _5685_/B _5292_/B _5703_/C _5398_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi221_1
X_7203_ _7404_/Q _7203_/A2 _7203_/B1 _7374_/Q _7208_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_99_641 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_7134_ _7938_/Q _7133_/S _7161_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_4346_ _7435_/Q _4347_/A2 _6622_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_99_685 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_113_495 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7065_ _7696_/Q _7194_/A2 _7194_/B1 _7664_/Q _7194_/C1 _7810_/Q _7068_/A2 VDD VSS
+ gf180mcu_fd_sc_mcu7t5v0__aoi222_1
Xclkbuf_leaf_75_csclk _7396_/CLK _7532_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
X_4277_ _7886_/Q _6520_/A1 _4527_/A1 _7373_/Q _4279_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_74_508 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6016_ hold512/Z _6021_/A2 _6017_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_2007 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_100_189 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_36_37 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_39_295 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_2018 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2029 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_82_563 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_27_446 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_7967_ _7967_/D _7320_/Z _4415_/A2 hold5/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XTAP_1339 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1328 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1317 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1306 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_427 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_168_602 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7898_ _7898_/D _7901_/RN _7898_/CLK _7898_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_70_747 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_23_641 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6918_ _7914_/Q _7913_/Q _6936_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_2
Xclkbuf_leaf_13_csclk _7592_/CLK _7901_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
X_6849_ _6849_/A1 _6767_/C _6849_/B1 _6849_/B2 _7433_/Q _6850_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi221_1
XFILLER_22_140 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_168_668 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_167_123 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_156_808 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_7_807 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_182_104 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_167_178 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_155_318 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_108_201 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_148_392 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xclkbuf_leaf_28_csclk _7825_/CLK _7853_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_108_256 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_163_373 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_123_215 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_151_579 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_117_40 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
Xhold380 _7858_/Q hold380/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
XFILLER_2_534 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_117_84 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_117_73 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xhold391 _7842_/Q hold391/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
XFILLER_104_495 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_77_357 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_58_571 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_46_744 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_61_703 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_45_221 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_73_574 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1851 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1840 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_60_224 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_1884 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1873 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1862 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_9_100 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_174_605 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_1895 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_41_482 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_146_318 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_9_144 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_115_705 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4200_ _7807_/Q _6350_/A1 _4569_/A1 _7392_/Q _4812_/A1 _7495_/Q _4201_/A2 VDD VSS
+ gf180mcu_fd_sc_mcu7t5v0__aoi222_1
X_5180_ _5648_/A1 _5774_/A1 _5752_/B1 _5066_/Z _5180_/C1 _5448_/A1 _5186_/A2 VDD VSS
+ gf180mcu_fd_sc_mcu7t5v0__aoi222_1
XFILLER_123_771 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4131_ hold118/Z _4217_/A2 _4893_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_95_154 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4062_ _7865_/Q _6469_/A1 _4219_/A2 input14/Z _4063_/A4 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_3_96 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_95_176 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_49_582 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_64_530 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7821_ _7821_/D _7901_/RN _7821_/CLK _7821_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_64_574 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_7752_ _7752_/D _7901_/RN _7755_/CLK _7752_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
X_4964_ _4965_/B _5363_/A2 _5774_/B2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_52_747 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3915_ _7683_/Q _6073_/A1 _6248_/A1 _7765_/Q _3916_/A4 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_6703_ _7661_/Q _6885_/A2 _6885_/B1 _7709_/Q _6705_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_32_460 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7683_ _7683_/D _7901_/RN _7821_/CLK _7683_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
X_4895_ _4448_/Z _4897_/A2 _4895_/B _7537_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_20_611 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_177_487 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_165_638 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3846_ hold124/Z hold118/Z _6090_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_4
XFILLER_20_666 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6634_ _6634_/A1 _7906_/Q _6661_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_4
X_6565_ _6565_/A1 _6565_/A2 _6565_/B _7903_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_3777_ input58/Z _3731_/Z _3777_/B1 _7964_/Q _3778_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_180_619 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5516_ _5648_/A1 _5608_/B _5176_/B _5690_/A1 _5530_/B _5517_/A4 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi221_1
X_6496_ hold41/Z _6502_/A2 _6496_/B _7874_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_160_321 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_145_384 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5447_ _5458_/C _5661_/A1 _5527_/A1 _5458_/B _5682_/A1 _5448_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai32_1
XFILLER_105_215 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_105_237 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_5378_ _5585_/A1 _5708_/A2 _5378_/B _5378_/C _5733_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi211_2
XFILLER_113_292 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_7117_ _7852_/Q _7193_/A2 _7193_/B1 _7634_/Q _7193_/C1 _7730_/Q _7121_/A1 VDD VSS
+ gf180mcu_fd_sc_mcu7t5v0__aoi222_1
XFILLER_101_432 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4329_ _7412_/Q _4329_/A2 _7334_/Q _4330_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_7048_ _7048_/A1 _7048_/A2 _7048_/A3 _7048_/A4 _7054_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand4_1
XFILLER_59_357 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_47_519 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_170_37 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_86_176 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_28_711 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_47_69 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_27_243 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_82_371 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1114 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1103 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1147 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1125 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1136 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1169 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1158 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_70_566 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_63_68 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_30_408 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_51_780 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_156_605 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_137_2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_128_318 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_10_132 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_155_115 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_10_176 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_155_159 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_163_181 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_151_354 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_78_600 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_909 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_120_730 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_104_270 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_92_135 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_92_179 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2371 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2360 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_33_235 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_34_747 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_34_758 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2393 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2382 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_61_555 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1692 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1681 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1670 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_3700_ _7703_/Q _3700_/ZN VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_159_465 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_147_627 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4680_ _7464_/Q hold55/Z _4680_/B hold69/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_147_649 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_147_638 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_146_126 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3631_ _7979_/Q _3735_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_174_479 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6350_ _6350_/A1 hold32/Z _6366_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_4
XFILLER_161_107 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5301_ _5301_/A1 _5303_/A4 _5301_/B _5359_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_155_682 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_6_670 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_52_2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_142_321 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6281_ hold90/Z _6281_/A2 _6281_/B _7773_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_5232_ _3722_/I _3723_/I _5006_/B _5006_/C _5303_/A4 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor4_4
XFILLER_130_527 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5163_ _5319_/C _5692_/B _5645_/A1 _5501_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor3_1
XFILLER_123_590 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_68_110 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_96_463 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_4114_ hold133/Z _3869_/I _4569_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_5094_ _5458_/B _5682_/A1 _5094_/B1 _5661_/A1 _5094_/C _5095_/C VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai221_1
XFILLER_111_785 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_96_496 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_84_636 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_69_699 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_68_176 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_56_316 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4045_ _7785_/Q _6299_/A1 hold119/I _7727_/Q _4249_/A2 input29/Z _4046_/A4 VDD VSS
+ gf180mcu_fd_sc_mcu7t5v0__aoi222_1
XFILLER_37_552 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_37_563 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_7804_ _7804_/D _7901_/RN _7805_/CLK _7804_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_64_382 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_25_747 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_219 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_208 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
X_5996_ hold73/Z _6004_/A2 _5996_/B hold385/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_24_246 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_25_769 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4947_ _4943_/Z _4956_/A2 _4979_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_2
X_7735_ _7735_/D _7961_/RN _7735_/CLK _7735_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_33_780 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_33_791 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_52_599 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_178_763 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_138_605 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7666_ _7666_/D _7901_/RN _7805_/CLK _7666_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
X_4878_ _4878_/A1 _7285_/A2 _4882_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_177_295 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3829_ hold630/I hold20/I _4275_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_4
XFILLER_20_474 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_20_463 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6617_ _7904_/Q _7905_/Q _6561_/Z _7435_/Q _6618_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai31_1
XFILLER_165_468 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7597_ _7597_/D _7961_/RN _7689_/CLK _7597_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_146_671 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6548_ hold525/Z _6553_/A2 _6549_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_161_641 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_145_181 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6479_ hold41/Z _6485_/A2 _6479_/B _7866_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_160_162 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_133_354 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xoutput260 _7571_/Q pll_bypass VDD VSS gf180mcu_fd_sc_mcu7t5v0__buf_8
Xoutput271 _7363_/Q pll_trim[0] VDD VSS gf180mcu_fd_sc_mcu7t5v0__buf_8
Xoutput293 _7369_/Q pll_trim[6] VDD VSS gf180mcu_fd_sc_mcu7t5v0__buf_8
Xoutput282 _7364_/Q pll_trim[1] VDD VSS gf180mcu_fd_sc_mcu7t5v0__buf_8
XFILLER_58_68 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_47_338 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_74_179 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_62_308 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_28_585 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_16_747 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_43_522 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_55_382 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_31_706 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_130_84 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_90_33 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_156_435 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_129_638 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_90_99 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_23_82 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_139_82 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_99_20 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_11_496 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_137_682 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_124_321 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_99_97 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_124_376 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_706 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_155_70 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_2_183 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_717 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_728 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_739 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_78_463 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_66_625 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_93_444 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_93_499 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_81_617 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_80_105 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_179_505 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_80_127 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_80_116 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5850_ hold692/Z _5851_/A2 _5851_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_34_566 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5781_ _5565_/Z _5781_/A2 _5782_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_1
XTAP_2190 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_4801_ _7487_/Q _4809_/S _4802_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_7520_ _7520_/D _7959_/RN _7958_/CLK _7520_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_4
X_4732_ _5903_/A2 hold32/Z _4742_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_2
X_7451_ hold4/Z _7901_/RN _7463_/CLK hold79/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_174_210 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_159_273 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_4663_ hold55/Z _4460_/Z _4664_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_9_73 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_30_772 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_175_777 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6402_ hold744/Z _6417_/A2 _6403_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_7382_ _7382_/D _7901_/RN _7810_/CLK _7382_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_128_671 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4594_ _4594_/A1 _7285_/A2 _4598_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_143_641 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_127_192 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6333_ _6333_/A1 _7285_/A2 _6349_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_4
XFILLER_170_460 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6264_ hold90/Z _6264_/A2 _6264_/B _7765_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_115_354 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5215_ _5200_/B _3727_/I _5421_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_142_195 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_8003_ _8003_/I _8003_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_6195_ hold722/Z _6208_/A2 _6196_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_5146_ _5643_/A2 _5752_/B1 _5186_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_97_783 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5077_ _5585_/A1 _5783_/A2 _5583_/C _5077_/C _5098_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi211_1
X_4028_ _7818_/Q hold134/I _6265_/A1 _7770_/Q hold108/I _8008_/I _4030_/A3 VDD VSS
+ gf180mcu_fd_sc_mcu7t5v0__aoi222_1
XFILLER_56_179 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_44_37 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_5979_ hold73/Z _5987_/A2 _5979_/B hold323/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_40_525 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_7718_ _7718_/D _7901_/RN _7799_/CLK _7718_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffsnq_1
XFILLER_100_54 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_40_569 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_178_582 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_166_744 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_21_783 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
Xclkbuf_1_1__f__1040_ clkbuf_0__1040_/Z _7226_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
X_7649_ _7649_/D _7961_/RN _7649_/CLK _7649_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_181_736 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_106_321 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_4_448 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_4_459 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_106_387 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_69_67 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_121_357 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_95_709 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_632 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_125_73 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_698 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_47_124 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_75_488 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_62_105 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_75_499 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_62_116 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_16_511 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_71_661 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_43_363 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_116_118 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_7_242 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_172_747 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_171_246 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_125_641 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_116_129 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
Xhold209 _7702_/Q hold209/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
XFILLER_7_286 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_152_460 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_124_151 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_98_536 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_525 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_514 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_503 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_5000_ _5600_/A1 _5363_/A2 _5658_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_4
XTAP_547 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_536 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_558 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_85_208 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_79_783 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_66_411 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_569 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_15_2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_27_809 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_38_124 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_38_179 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_81_447 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_81_425 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_53_138 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6951_ _6955_/A4 _6951_/A2 _7188_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_4
X_5902_ hold90/Z _5902_/A2 _5902_/B _7595_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_6882_ _7757_/Q _6882_/A2 _6882_/B1 _7495_/Q _6888_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_179_335 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_61_160 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5833_ _7565_/Q _5840_/A2 _5834_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_50_812 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_179_357 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_14_29 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_148_733 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_5764_ _5579_/B _5764_/A2 _5744_/Z _5746_/Z _5805_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor4_2
X_7503_ _7503_/D _7912_/CLK _7503_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_4715_ _7443_/Q _4718_/A1 _4718_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_5695_ _5706_/A2 _5625_/Z _5725_/A2 _5691_/Z _5695_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__and4_1
X_4646_ _3830_/Z hold68/Z _4647_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_107_107 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7434_ _7434_/D _7961_/RN _7940_/CLK _7434_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_2
Xhold721 _7701_/Q hold721/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
X_7365_ _7365_/D _7961_/RN _7565_/CLK _7365_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffsnq_2
Xhold710 _7504_/Q hold710/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
X_4577_ hold616/Z _4578_/A2 _4578_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_162_257 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
Xhold754 _3803_/Z hold754/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
X_6316_ _6316_/A1 _7285_/A2 _6332_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_4
Xhold732 _7862_/Q hold732/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
Xhold743 _7620_/Q hold743/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
XFILLER_171_780 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7296_ _7901_/RN _4334_/Z _7296_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_131_611 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_116_696 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
Xhold765 _7870_/Q hold765/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
XFILLER_130_143 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_115_195 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_103_357 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_77_709 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6247_ _4454_/Z _6247_/A2 _6247_/B _7757_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_6178_ hold568/Z _6191_/A2 _6179_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_85_720 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5129_ _5705_/A2 _5179_/B _5657_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_84_230 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_55_69 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_57_499 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_111_31 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_111_20 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_40_311 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_41_812 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_13_558 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_154_725 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_138_276 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_126_405 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_154_747 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_107_641 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_134_460 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_106_162 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_136_83 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_136_94 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_96_21 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_121_154 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_67_208 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_48_400 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_484 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xhold81 hold81/I hold81/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
Xhold92 hold92/I hold92/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
Xhold70 hold70/I hold70/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
XFILLER_91_712 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_48_477 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_152_93 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_35_138 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_90_277 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_32_812 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_50_108 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_31_377 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_176_349 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_129_232 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_129_221 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5480_ _5538_/A1 _5026_/Z _5480_/A3 _5652_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand3_1
X_4500_ hold47/Z _4504_/A2 _4500_/B hold541/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_172_522 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_6_52 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4431_ input1/Z input36/Z _4431_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_160_717 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_132_408 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_99_812 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7150_ _7853_/Q _7193_/A2 _7189_/A2 _7715_/Q _7153_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_4362_ _6623_/B _4362_/A2 _7435_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_4293_ _4309_/S _4300_/C VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_6101_ hold426/Z _6106_/A2 _6102_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_112_132 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_112_110 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7081_ _7935_/Q _7133_/S _7082_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_59_709 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_140_485 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_140_463 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_100_316 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_98_377 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6032_ hold41/Z _6038_/A2 _6032_/B hold443/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
XTAP_366 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_39_411 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_79_580 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_377 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_399 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_388 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_26_105 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_39_499 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7983_ _7983_/I _7983_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XPHY_28 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_17 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
X_6934_ _7912_/Q _7911_/Q _6941_/A2 _6908_/Z _7201_/B1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor4_4
XPHY_39 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_23_812 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_179_132 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_62_491 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_6865_ _7756_/Q _6882_/A2 _6894_/C1 _7403_/Q _6865_/C _6867_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi221_1
X_6796_ _7763_/Q _6892_/A2 _6892_/B1 _7729_/Q _6799_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_5816_ _4454_/Z _5816_/A2 _5816_/B hold707/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_148_530 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5747_ _5747_/A1 _5747_/A2 _5756_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_22_388 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_108_416 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5678_ _5678_/A1 _5064_/B _5678_/A3 _5679_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor3_1
XFILLER_136_747 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7417_ hold81/Z _7901_/RN _7461_/CLK _7991_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
X_4629_ _7992_/I _4652_/A1 _4632_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_135_246 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_173_26 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
Xhold562 _7456_/Q hold562/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
XFILLER_150_205 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_116_460 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xhold551 _7367_/Q hold551/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
Xhold540 hold540/I _4500_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
XFILLER_1_215 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_7348_ _7348_/D _7961_/RN _7353_/CLK _7348_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffsnq_2
X_7279_ _7279_/A1 _7279_/A2 _7279_/B _7517_/Q _7958_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi211_1
Xhold584 _7661_/Q hold584/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
Xclkbuf_3_5__f_csclk clkbuf_0_csclk/Z _7825_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_89_344 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
Xhold573 _7530_/Q hold573/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
Xhold595 _7469_/Q hold595/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
XFILLER_104_699 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_131_496 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_58_742 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_181_4 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_85_550 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_73_712 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_17_105 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_45_425 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_167_2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_45_469 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_82_34 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_73_789 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_72_277 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_14_812 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_32_108 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_9_304 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_40_152 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_41_653 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_154_522 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_126_213 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_5_521 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_154_599 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_135_780 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_107_460 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_99_119 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_122_463 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_122_474 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_68_506 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_1_771 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_163_70 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_83_509 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_64_701 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
Xinput160 wb_rstn_i _7959_/RN VDD VSS gf180mcu_fd_sc_mcu7t5v0__buf_12
XFILLER_76_583 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_63_211 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_48_285 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_91_531 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_64_756 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_36_458 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4980_ _5741_/A1 _4993_/B _5735_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_4
XFILLER_17_661 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_51_428 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3931_ _7674_/Q _6056_/A1 _5920_/A1 _7610_/Q hold134/I _7820_/Q _3955_/A2 VDD VSS
+ gf180mcu_fd_sc_mcu7t5v0__aoi222_4
XFILLER_177_636 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_149_316 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3862_ hold123/Z _3787_/Z hold127/Z _3794_/Z _4151_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand4_4
X_6650_ _6878_/A2 _6664_/A3 _6662_/A3 _6894_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor3_4
X_5601_ _5783_/A2 _5668_/A2 _5668_/C _5612_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_82_2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6581_ _6586_/A1 _6581_/A2 _6663_/A4 _6586_/B _7907_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand4_1
XFILLER_176_179 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3793_ hold153/Z input58/Z _7414_/Q _3793_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_5532_ _5648_/A2 _5179_/B _5555_/B _5555_/C _5743_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XFILLER_145_511 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_118_747 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_145_577 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_145_566 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5463_ _5643_/A2 _5783_/A2 _5585_/B _5772_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi21_1
Xclkbuf_leaf_9_csclk clkbuf_leaf_9_csclk/I _7897_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_8_392 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5394_ _5394_/A1 _5709_/A2 _5394_/B _5415_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_160_514 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4414_ _7919_/Q _7576_/Q _7580_/Q _4414_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_7202_ _7408_/Q _7202_/A2 _7202_/B1 _7398_/Q _7386_/Q _7202_/C2 _7208_/A1 VDD VSS
+ gf180mcu_fd_sc_mcu7t5v0__aoi222_1
XFILLER_132_238 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7133_ _7133_/I0 _7937_/Q _7133_/S _7937_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_4345_ _7904_/Q _7905_/Q _4347_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_141_783 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_98_174 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_143_29 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_101_658 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_100_102 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_7064_ _7850_/Q _7193_/A2 _7193_/B1 _7632_/Q _7193_/C1 _7728_/Q _7068_/A1 VDD VSS
+ gf180mcu_fd_sc_mcu7t5v0__aoi222_1
X_4276_ input52/Z _5886_/A1 _4888_/A1 _7535_/Q _4279_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_6015_ hold41/Z _6021_/A2 _6015_/B hold518/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_39_241 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_39_230 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_100_179 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_67_572 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_55_712 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_2019 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2008 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_82_531 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7966_ _7966_/D _7319_/Z _4415_/A2 hold1/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XTAP_1329 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1318 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1307 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_14_108 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_7897_ _7897_/D _7901_/RN _7897_/CLK _7897_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffsnq_1
X_6917_ _6953_/A2 _6955_/A4 _6908_/Z _7207_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor3_4
X_6848_ _6848_/A1 _6848_/A2 _6848_/A3 _6849_/B2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor3_1
XFILLER_23_653 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_52_37 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_168_37 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6779_ _7433_/Q _7924_/Q _6779_/B _6781_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_10_347 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_182_138 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_136_522 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_109_736 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_6_318 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_151_503 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_117_780 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_117_30 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_117_63 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_117_52 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xhold370 _7882_/Q hold370/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
Xhold381 _7576_/Q hold381/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
XFILLER_104_463 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_89_141 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xhold392 _7834_/Q hold392/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
XFILLER_77_89 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_58_550 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_133_73 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_92_328 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_93_66 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_46_756 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_73_586 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_33_406 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_33_428 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1852 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1841 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1830 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_61_759 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_158_102 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1885 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1874 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1863 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_13_141 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_158_146 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1896 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_158_179 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_42_70 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_182_661 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_182_650 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_182_694 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_182_683 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_170_812 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_154_374 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_5_373 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_154_396 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_123_783 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4130_ hold133/Z _3881_/Z _4609_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_122_282 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_95_144 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4061_ input46/Z _4275_/A2 _5817_/A1 _7561_/Q _6282_/A1 _7777_/Q _4063_/A3 VDD VSS
+ gf180mcu_fd_sc_mcu7t5v0__aoi222_1
XFILLER_37_734 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_37_723 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_37_712 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7820_ _7820_/D _7901_/RN _7820_/CLK _7820_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_64_542 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_91_361 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_64_586 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_52_726 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4963_ _5069_/A2 _4930_/Z _4953_/Z _4963_/A4 _5363_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand4_4
X_7751_ _7751_/D _7901_/RN _7753_/CLK _7751_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
X_7682_ _7682_/D _7901_/RN _7698_/CLK _7682_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
X_3914_ _7731_/Q hold119/I _6384_/A1 _7829_/Q _3916_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_6702_ _6702_/A1 _6702_/A2 _6702_/A3 _6706_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_177_433 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_149_124 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_4894_ hold658/Z _4897_/A2 _4895_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_6633_ _7907_/Q _6633_/A2 _6665_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_164_105 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3845_ _3835_/Z hold113/Z _6209_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_4
XFILLER_20_656 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_177_499 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_164_127 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_138_29 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6564_ _7435_/Q _6569_/A3 _6564_/B _7902_/Q _6565_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai211_1
X_3776_ _7411_/Q _3730_/Z _4380_/A2 _3777_/B1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand3_1
X_5515_ _5179_/B _5672_/A2 _5550_/B _5517_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_6495_ hold358/Z _6502_/A2 _6496_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_161_812 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_145_363 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5446_ _5446_/A1 _5446_/A2 _5446_/A3 _5520_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_106_739 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_160_344 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_133_547 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_121_709 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5377_ _5378_/B _5711_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_7116_ _7116_/A1 _7116_/A2 _7116_/A3 _7116_/A4 _7130_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand4_1
X_4328_ _7415_/Q _3734_/Z _4329_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_7047_ _7655_/Q _7189_/C1 _7207_/B1 _7719_/Q _7048_/A4 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_4259_ _7660_/Q _6039_/A1 _5855_/A1 _7982_/I _4260_/A4 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_101_499 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_27_211 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_103_65 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1104 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_7949_ _7949_/D _7949_/CLK _7949_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_70_534 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_1137 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1115 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1126 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_15_428 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_27_299 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_168_400 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1159 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1148 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_247 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_42_258 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_50_291 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_7_638 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_170_108 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_152_812 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_136_396 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_128_84 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_128_95 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_88_33 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_2_321 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_111_208 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_105_783 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_104_282 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_77_144 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_77_133 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_19_701 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_19_712 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_46_531 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_19_778 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_179_709 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2350 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2361 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_160_93 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_73_394 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_46_597 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2394 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2383 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2372 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1660 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_61_578 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_61_567 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1693 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1682 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1671 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
Xclkbuf_leaf_74_csclk _7396_/CLK _7625_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_159_499 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_159_488 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_146_116 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3630_ _7980_/Q _4424_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_5300_ _5166_/C _5300_/A2 _5360_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_143_812 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_127_352 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6280_ hold471/Z _6281_/A2 _6281_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
Xclkbuf_leaf_89_csclk _7396_/CLK _7570_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
X_5231_ _4915_/Z _5303_/A3 _5258_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_103_709 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_45_2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5162_ _5218_/B _5498_/B _5162_/B _5162_/C _5187_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_69_645 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5093_ _5087_/C _4898_/Z _5424_/A1 _5094_/C VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand3_1
Xclkbuf_leaf_12_csclk _7592_/CLK _7900_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
X_4113_ hold20/Z hold118/Z _4878_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_69_689 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_4044_ _7687_/Q _6090_/A1 _6073_/A1 _7679_/Q _6141_/A1 _7711_/Q _4046_/A3 VDD VSS
+ gf180mcu_fd_sc_mcu7t5v0__aoi222_1
XFILLER_17_29 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_49_380 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_49_391 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
Xclkbuf_leaf_27_csclk _7592_/CLK _7877_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
X_7803_ _7803_/D _7901_/RN _7819_/CLK _7803_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_52_534 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7734_ _7734_/D _7901_/RN _7818_/CLK _7734_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffsnq_1
XPHY_209 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
X_5995_ hold384/Z _6004_/A2 _5996_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_40_707 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4946_ _4946_/A1 _5230_/A1 _4917_/Z _5369_/B _4955_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai22_2
XFILLER_33_770 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7665_ _7665_/D _7901_/RN _7820_/CLK _7665_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_177_263 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4877_ _4454_/Z _4877_/A2 _4877_/B _7530_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_165_425 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3828_ hold20/Z _4620_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_7596_ _7596_/D _7961_/RN _7689_/CLK _7596_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
X_6616_ _7916_/Q _6611_/B _6616_/B _7916_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_6547_ hold41/Z _6553_/A2 _6547_/B _7898_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_152_108 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_134_812 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3759_ _4292_/B _3759_/A2 _7974_/Q _3760_/B2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_161_631 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_145_193 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_6478_ hold500/Z _6485_/A2 _6479_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_160_130 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_133_366 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_5429_ _5624_/A1 _5648_/B2 _5685_/B _5614_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
Xoutput261 _7557_/Q pll_dco_ena VDD VSS gf180mcu_fd_sc_mcu7t5v0__buf_8
Xoutput250 _4435_/Z pad_flash_csb_oe VDD VSS gf180mcu_fd_sc_mcu7t5v0__buf_8
XFILLER_160_196 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xoutput294 _7370_/Q pll_trim[7] VDD VSS gf180mcu_fd_sc_mcu7t5v0__buf_8
Xoutput272 _7357_/Q pll_trim[10] VDD VSS gf180mcu_fd_sc_mcu7t5v0__buf_8
Xoutput283 _7351_/Q pll_trim[20] VDD VSS gf180mcu_fd_sc_mcu7t5v0__buf_8
XFILLER_59_144 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_87_475 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_101_296 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_28_531 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_28_520 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_130_30 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_43_567 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_129_628 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_128_105 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_144_609 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_128_149 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_128_138 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_171_428 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_125_812 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_99_54 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_136_193 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_151_141 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_151_152 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_3_641 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_707 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_151_185 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_97_217 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_718 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_729 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_38_328 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_48_91 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_76 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_34_534 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2180 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_4800_ _7219_/A1 _4809_/S _4800_/B _7486_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
XTAP_2191 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_5780_ _5372_/Z _5780_/A2 _5780_/B _5781_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_21_228 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_175_712 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_1490 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_4731_ hold47/Z _4731_/A2 _4731_/B _7449_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_7450_ hold17/Z _7901_/RN _7450_/CLK _7450_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
X_4662_ _7983_/I _4685_/A1 _4665_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_147_425 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6401_ _6401_/A1 _7285_/A2 _6417_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_4
X_7381_ _7381_/D _7901_/RN _7746_/CLK _7381_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_134_108 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_116_812 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4593_ _4454_/Z _4593_/A2 _4593_/B _7400_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_143_631 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6332_ hold90/Z _6332_/A2 _6332_/B _7797_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_115_311 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6263_ hold375/Z _6264_/A2 _6264_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_115_366 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_88_206 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_170_472 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5214_ _5669_/A1 _5087_/B _5218_/C VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_142_163 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_8002_ _8002_/I _8002_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_6194_ _4448_/Z _6208_/A2 _6194_/B _7732_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_5145_ _5643_/A2 _5608_/B _5739_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_96_250 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_57_615 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5076_ _5669_/B _4996_/Z _5465_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_4027_ _7744_/Q _6209_/A1 _6248_/A1 _7762_/Q _4030_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_72_618 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_13_707 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_25_567 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5978_ hold322/Z _5987_/A2 _5979_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_80_673 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_13_718 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4929_ _5195_/B _4914_/Z _5210_/A3 _4951_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor3_2
X_7717_ _7717_/D _7901_/RN _7799_/CLK _7717_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffsnq_1
XFILLER_100_44 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_100_88 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_60_37 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_20_250 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_7648_ _7648_/D _7961_/RN _7648_/CLK _7648_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_176_37 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_165_244 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_121_6 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_20_272 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_153_428 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_119_650 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_107_812 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7579_ _7579_/D _7961_/RN _7580_/CLK _7579_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_180_247 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_109_42 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_133_141 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_122_804 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_79_239 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_88_784 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_85_23 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_87_294 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_87_283 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_85_67 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_48_659 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_90_404 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_141_73 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_90_426 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_90_415 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_16_534 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_28_372 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_90_459 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_70_183 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_157_712 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_156_211 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_117_609 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_11_283 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_8_733 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_7_221 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_116_108 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_125_631 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_152_483 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_152_472 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_515 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_504 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_140_656 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_124_196 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_548 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_537 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_526 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_78_250 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_559 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_38_103 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_39_637 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_39_648 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6950_ _6950_/A1 _6950_/A2 _6955_/A4 _7204_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor3_4
XFILLER_54_607 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_54_618 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_93_286 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5901_ hold300/Z _5902_/A2 _5902_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_53_106 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_81_459 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6881_ _7530_/Q _6881_/A2 _6881_/B1 _7524_/Q _6888_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_179_325 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_62_673 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5832_ _4454_/Z _5840_/A2 _5832_/B _7564_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_5763_ _5763_/A1 _5698_/B _5763_/A3 _5763_/A4 _5792_/B1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor4_2
X_4714_ _4718_/A1 hold86/Z _4714_/B hold87/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_7502_ _7502_/D _7912_/CLK _7502_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_148_756 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5694_ _5424_/Z _5763_/A1 _5723_/A1 _5694_/A4 _5696_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor4_1
XFILLER_175_586 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4645_ hold197/Z _4652_/A1 _4648_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_135_428 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_30_29 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_7433_ _7433_/D _7961_/RN _7940_/CLK _7433_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_4
XFILLER_162_247 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_146_29 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_135_439 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7364_ _7364_/D _7961_/RN _7565_/CLK _7364_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffsnq_1
Xhold700 hold700/I _7356_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
X_4576_ _4448_/Z _4578_/A2 _4576_/B _7393_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
Xhold711 _7409_/Q hold711/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
XFILLER_143_450 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_115_141 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6315_ hold90/Z _6315_/A2 _6315_/B _7789_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
Xhold744 _7830_/Q hold744/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
Xhold733 _7838_/Q hold733/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
Xhold755 hold755/I _7571_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
Xhold722 _7733_/Q hold722/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
X_7295_ _7901_/RN _4334_/Z _7295_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_116_686 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_115_185 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_115_152 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_103_303 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xhold766 _7814_/Q hold766/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
X_6246_ hold570/Z _6247_/A2 _6247_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_6177_ _4448_/Z _6191_/A2 _6177_/B _7724_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_97_570 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_39_49 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5128_ _5600_/A1 _5797_/B _5527_/A1 _5166_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor3_1
XFILLER_69_283 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_57_478 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5059_ _5195_/B _5016_/B _5692_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_4
XFILLER_84_275 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_72_459 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_41_802 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_139_712 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_138_211 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_71_69 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_166_531 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_139_767 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_21_570 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_181_512 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_153_203 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_139_778 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_138_266 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_138_255 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_119_491 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_119_480 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_112_2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_181_567 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_153_269 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_136_62 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_121_100 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_106_174 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_122_656 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_122_678 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_121_144 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_95_507 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xhold82 hold82/I hold82/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
Xhold71 hold71/I hold71/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
Xhold60 hold60/I hold60/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
XFILLER_152_72 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_29_93 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_48_456 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xhold93 hold93/I hold93/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
XFILLER_75_297 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_75_286 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_45_70 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_44_673 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_31_334 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_31_345 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_31_367 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_129_277 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_172_534 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_145_737 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_117_428 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4430_ _4396_/S input63/Z _4430_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_144_247 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_6_64 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_98_323 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6100_ hold41/Z _6106_/A2 _6100_/B _7688_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_4361_ _7433_/Q _4361_/A2 _4361_/A3 _4362_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand3_1
X_7080_ _7433_/Q _7934_/Q _7078_/Z _7080_/B2 _7082_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_4292_ _7414_/Q _4292_/A2 _4292_/B _4309_/S VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_4
XFILLER_98_389 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_79_570 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6031_ hold442/Z _6038_/A2 _6032_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_367 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_389 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_378 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_39_478 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_82_724 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_7982_ _7982_/I _7982_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XPHY_18 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_29 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
X_6933_ _6941_/A2 _6951_/A2 _7193_/B1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_4
XFILLER_34_161 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6864_ _6864_/A1 _6864_/A2 _6864_/A3 _6865_/C VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_179_144 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_90_790 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_62_481 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5815_ hold705/Z _5816_/A2 hold706/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_22_312 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6795_ _7827_/Q _6891_/A2 _6891_/B1 _7673_/Q _6891_/C1 _7779_/Q _6799_/A1 VDD VSS
+ gf180mcu_fd_sc_mcu7t5v0__aoi222_1
XFILLER_50_676 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_179_199 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5746_ _5380_/I _5501_/Z _5524_/I _5746_/A4 _5746_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__or4_1
XFILLER_22_378 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5677_ hold18/I _5520_/C _5677_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__and2_1
X_4628_ _4652_/A1 hold80/Z _4628_/B hold81/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_148_597 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_136_737 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_7416_ _7416_/D _7901_/RN _7450_/CLK _7990_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_163_567 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_151_707 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
Xhold530 _7777_/Q hold530/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
Xhold563 _4740_/Z _7456_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
Xhold552 hold552/I _4515_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
Xhold541 hold541/I _7360_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
XFILLER_2_717 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_4559_ _4559_/A1 _7285_/A2 _4563_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_7347_ _7347_/D _7961_/RN _7353_/CLK _7347_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffsnq_1
X_7278_ _7278_/A1 _7277_/B _7278_/B _7957_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi21_1
Xhold585 hold585/I _6043_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
Xhold596 _7477_/Q hold596/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
Xhold574 _7402_/Q hold574/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
X_6229_ hold567/Z _6242_/A2 _6230_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_106_43 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_103_144 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_77_529 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_103_177 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_890 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_57_286 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_122_64 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_73_779 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_45_448 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_72_256 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_26_673 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_25_161 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_158_328 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_15_73 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_40_175 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_41_698 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_139_564 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_154_534 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_127_737 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_126_203 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_147_61 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_126_247 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_147_94 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_99_109 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_5_566 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_68_518 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_1_761 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_110_626 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_282 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_1_783 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
Xinput161 wb_sel_i[0] _7236_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
Xinput150 wb_dat_i[2] _7252_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_76_551 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_48_242 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_76_595 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_49_787 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_49_798 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_63_223 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3930_ _7884_/Q _6503_/A1 hold26/I _3927_/Z _6005_/A1 _7650_/Q _3955_/A1 VDD VSS
+ gf180mcu_fd_sc_mcu7t5v0__aoi222_4
XFILLER_51_407 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_176_103 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3861_ _3817_/I hold118/Z hold119/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_4
XFILLER_32_676 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3792_ _7506_/Q hold104/Z _3792_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__and2_1
X_5600_ _5600_/A1 _5797_/B _4993_/C _5458_/B _5600_/B2 _5668_/C VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai32_1
X_6580_ _7432_/Q _4352_/B _6586_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_2
X_5531_ _5543_/B _5539_/A3 _5541_/A4 _5555_/C VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor3_1
XFILLER_75_2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_117_225 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_172_342 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5462_ _4969_/C _5604_/A2 _5658_/B _5608_/B _5462_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__or4_1
X_7201_ _7372_/Q _7201_/A2 _7201_/B1 _7508_/Q _7206_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_160_526 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_160_504 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5393_ _5380_/I _5565_/A2 _5581_/C _5394_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__or3_1
XFILLER_132_228 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_126_770 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4413_ _7917_/Q _7577_/Q _7580_/Q _4413_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_4344_ _4344_/I _7520_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_7132_ _7433_/Q _7132_/A2 _7132_/B _7133_/I0 VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_140_250 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7063_ _7063_/A1 _7063_/A2 _7063_/A3 _7063_/A4 _7078_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand4_1
XFILLER_59_507 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_141_795 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_140_272 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4275_ input43/Z _4275_/A2 _4549_/A1 _7383_/Q _4279_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_6014_ hold517/Z _6021_/A2 _6015_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_55_702 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_39_286 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2009 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_94_392 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1319 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1308 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_82_587 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_7965_ _7965_/D _7318_/Z _7977_/CLK _7965_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_54_256 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7896_ _7896_/D _7901_/RN _7900_/CLK _7896_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_23_621 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6916_ _6950_/A1 _6941_/A2 _6908_/Z _7189_/B1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor3_4
X_6847_ _6847_/A1 _6847_/A2 _6847_/A3 _6848_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand3_1
X_6778_ _7079_/A1 _6767_/C _6778_/B _7433_/Q _6779_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi211_1
X_5729_ _5791_/A2 _5761_/A2 _5762_/A4 _5730_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_176_692 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_148_383 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_136_534 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_108_247 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_117_42 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xhold371 _7890_/Q hold371/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
Xhold360 hold360/I _7625_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
XFILLER_132_762 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_132_751 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
Xhold393 _7674_/Q hold393/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
Xhold382 _7658_/Q hold382/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
XFILLER_78_805 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_131_283 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_92_318 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_85_381 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_73_554 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_45_212 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_33_418 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_45_278 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1842 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1831 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1820 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_61_749 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_14_621 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1875 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1864 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1853 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1897 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1886 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_14_676 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_139_350 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_41_495 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_9_168 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_127_567 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_181_161 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_181_194 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_122_250 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_96_602 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_110_456 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_110_445 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4060_ _7615_/Q _5937_/A1 _6226_/A1 _7751_/Q _4063_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_110_489 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_67_90 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_76_392 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7750_ _7750_/D _7901_/RN _7755_/CLK _7750_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffsnq_1
X_4962_ _5369_/B _4943_/Z _5603_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_4
XFILLER_91_373 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_64_598 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_24_429 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_51_215 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_149_103 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3913_ _7715_/Q _6141_/A1 _6265_/A1 _7773_/Q _3916_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_7681_ _7681_/D _7901_/RN _7691_/CLK _7681_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
X_6701_ _7376_/Q _6882_/A2 _6880_/A2 _7815_/Q _6702_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_4893_ _4893_/A1 _7285_/A2 _4897_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_3844_ _4212_/A2 _4075_/B _4488_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_4
XFILLER_20_602 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6632_ _7910_/Q _6664_/A3 _6662_/A3 _6881_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor3_4
XFILLER_22_19 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_164_139 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_158_670 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6563_ _6563_/I _6565_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_3775_ _7965_/Q _3738_/Z _4380_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_5514_ _5514_/A1 _5514_/A2 _5514_/A3 _5514_/A4 _5518_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand4_1
XFILLER_118_534 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6494_ hold73/Z _6502_/A2 _6494_/B _7873_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_5445_ _5783_/B _5757_/B _5445_/A3 _5445_/A4 _5446_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor4_1
XFILLER_172_172 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5376_ _5371_/C _5392_/B2 _5376_/B _5378_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_114_751 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7115_ _7690_/Q _7189_/B1 _7189_/C1 _7658_/Q _7115_/C _7116_/A4 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi221_1
XFILLER_141_570 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_113_283 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_99_473 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4327_ _7964_/Q _7335_/Q _4327_/S _7335_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_7046_ _7727_/Q _7193_/C1 _7196_/B1 _7639_/Q _7048_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_4258_ _7716_/Q _6158_/A1 _4878_/A1 _7531_/Q _4260_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_86_189 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_74_318 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4189_ input72/Z _5903_/A1 _4232_/A2 input35/Z _4584_/A1 _7398_/Q _4203_/A3 VDD VSS
+ gf180mcu_fd_sc_mcu7t5v0__aoi222_2
XFILLER_55_521 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_103_55 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1105 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_55_565 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_103_99 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_7948_ _7948_/D _7949_/CLK _7948_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_70_524 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_1138 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1116 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1127 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1149 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_7879_ _7879_/D input75/Z _7887_/CLK _7879_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffsnq_1
XFILLER_155_117 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_6_105 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_109_567 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_164_673 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_163_161 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_151_301 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_3_812 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_136_386 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_78_602 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_5_2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_132_592 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_120_721 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_104_272 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_104_250 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
Xhold190 hold190/I _7888_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
XFILLER_78_613 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_78_624 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_78_635 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_66_808 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_93_638 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_58_392 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xclkbuf_leaf_8_csclk clkbuf_leaf_9_csclk/I _7898_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_73_351 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_18_256 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_18_245 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_46_565 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2351 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2362 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2340 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_33_215 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_34_727 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_34_749 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_34_738 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2395 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2384 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2373 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_159_401 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_1650 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_61_557 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1694 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1683 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1672 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1661 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_53_81 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_53_70 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_174_404 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_169_70 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_53_92 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_174_459 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_146_139 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_182_492 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_170_621 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_154_172 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5230_ _5230_/A1 _5054_/Z _5685_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_4
XFILLER_5_171 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_170_676 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_69_602 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5161_ _3723_/I _5579_/B _5162_/C VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_142_389 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_123_570 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_111_732 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_111_721 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_38_2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5092_ _5058_/Z _5456_/A2 _5114_/A3 _5776_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand3_2
XFILLER_110_242 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_84_605 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4112_ hold133/Z hold156/Z _4614_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_84_638 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4043_ _7735_/Q _6192_/A1 _6124_/A1 _7703_/Q _6107_/A1 _7695_/Q _4046_/A2 VDD VSS
+ gf180mcu_fd_sc_mcu7t5v0__aoi222_1
XFILLER_56_318 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7802_ _7802_/D _7901_/RN _7802_/CLK _7802_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
X_5994_ _4460_/Z _6004_/A2 _5994_/B hold177/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_4945_ _4900_/Z _4915_/Z _4945_/B1 _5022_/B _4956_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_2
X_7733_ _7733_/D _7961_/RN _7733_/CLK _7733_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffsnq_1
XFILLER_149_29 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7664_ _7664_/D _7901_/RN _7851_/CLK _7664_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
X_4876_ hold573/Z _4877_/A2 _4877_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_177_286 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3827_ hold19/Z _3925_/A2 _3790_/Z _3794_/Z hold20/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand4_4
X_7595_ _7595_/D input75/Z _7865_/CLK _8005_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_20_476 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_20_454 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6615_ _7916_/Q _6586_/B _6611_/B _6616_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_137_139 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6546_ hold379/Z _6553_/A2 _6547_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_3758_ _7975_/Q _3765_/A1 _3759_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_146_673 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_146_662 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_145_161 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_145_150 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_161_621 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_3689_ _7785_/Q _3689_/ZN VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_6477_ hold73/Z _6485_/A2 _6477_/B _7865_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_5428_ _5482_/B2 _5510_/A2 _5793_/B _5789_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi21_1
Xoutput251 _4423_/Z pad_flash_io0_do VDD VSS gf180mcu_fd_sc_mcu7t5v0__buf_8
XFILLER_0_804 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xoutput262 _7558_/Q pll_div[0] VDD VSS gf180mcu_fd_sc_mcu7t5v0__buf_8
Xoutput240 _7984_/Z mgmt_gpio_out[3] VDD VSS gf180mcu_fd_sc_mcu7t5v0__buf_8
X_5359_ _5359_/A1 _5359_/A2 _5636_/A1 _5359_/B _5360_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai31_1
XFILLER_114_581 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
Xoutput273 _7358_/Q pll_trim[11] VDD VSS gf180mcu_fd_sc_mcu7t5v0__buf_8
Xoutput295 _7355_/Q pll_trim[8] VDD VSS gf180mcu_fd_sc_mcu7t5v0__buf_8
Xoutput284 _7352_/Q pll_trim[21] VDD VSS gf180mcu_fd_sc_mcu7t5v0__buf_8
XFILLER_58_37 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_114_592 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_99_292 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_87_443 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_59_134 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_75_638 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_74_104 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7029_ _7933_/Q _7133_/S _7030_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_101_286 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_74_126 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_28_510 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_114_98 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_28_543 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_70_321 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_15_215 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_16_738 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_130_53 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_70_354 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_24_782 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_30_207 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_142_2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_129_618 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_23_73 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_156_459 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_139_73 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_7_425 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_125_802 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_152_676 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_3_631 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_152_687 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_124_389 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_105_570 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_708 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_719 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_66_605 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_38_318 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_65_137 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_80_118 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2170 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_61_354 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2192 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2181 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1491 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1480 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_4730_ hold350/Z _4731_/A2 _4731_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_174_212 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_159_286 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_4661_ _4685_/A1 hold37/Z _4661_/B hold38/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_147_415 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7380_ _7380_/D _7901_/RN _7746_/CLK _7380_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
X_6400_ hold90/Z _6400_/A2 _6400_/B _7829_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_80_90 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6331_ hold387/Z _6332_/A2 _6332_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_128_673 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4592_ hold575/Z _4593_/A2 _4593_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_170_451 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_142_131 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_142_120 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6262_ hold68/Z _6264_/A2 _6262_/B _7764_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_5213_ _4906_/Z _5373_/A3 _5373_/A4 _5405_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand3_4
XFILLER_142_175 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8001_ _8001_/I _8001_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_6193_ hold769/Z _6208_/A2 _6194_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_5144_ _5543_/C _5689_/A2 _5543_/B _5499_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor3_1
XFILLER_69_443 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_97_796 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_28_29 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5075_ _5603_/A1 _4993_/B _5663_/A1 _5583_/C VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor3_2
XFILLER_84_479 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4026_ _7826_/Q _6384_/A1 _5828_/A1 _7567_/Q _6537_/A1 _7898_/Q _4030_/A1 VDD VSS
+ gf180mcu_fd_sc_mcu7t5v0__aoi222_1
XFILLER_25_513 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_53_811 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_52_321 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5977_ _4460_/Z _5987_/A2 _5977_/B hold250/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_178_540 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_4928_ _4914_/Z _5210_/A3 _5195_/B _5069_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_4
X_7716_ _7716_/D _7901_/RN _7805_/CLK _7716_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffsnq_1
XFILLER_100_34 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_165_212 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_100_67 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_20_240 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_7647_ _7647_/D _7961_/RN _7692_/CLK _7647_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_138_459 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_20_262 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4859_ hold752/Z _4862_/A2 _4860_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_118_150 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_109_32 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_4_406 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7578_ _7578_/D _7961_/RN _7580_/CLK _7578_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_134_621 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_119_695 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_106_312 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6529_ hold371/Z _6536_/A2 _6530_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_134_676 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_106_345 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_69_36 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_161_495 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_106_389 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_102_551 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_667 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_48_605 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_75_446 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
Xclkbuf_leaf_73_csclk _7396_/CLK _7642_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_85_79 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_56_660 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_141_41 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_18_84 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_71_641 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xclkbuf_leaf_88_csclk _7396_/CLK _7353_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_43_332 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_43_354 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_169_540 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_156_201 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
Xclkbuf_leaf_11_csclk _7592_/CLK _7899_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_12_763 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_156_278 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_171_215 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_171_248 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xclkbuf_leaf_26_csclk _7825_/CLK _7844_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_140_602 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_125_698 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_124_175 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_516 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_505 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_549 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_538 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_527 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_3_494 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_79_785 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_79_763 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_39_605 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_120_392 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_94_744 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_78_295 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_66_413 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_38_126 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_94_788 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_93_232 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5900_ hold68/Z _5902_/A2 _5900_/B _7594_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_81_438 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_19_351 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_34_310 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_34_321 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_6880_ _7961_/Q _6880_/A2 _6880_/B1 _7410_/Q _7477_/Q _6880_/C2 _6888_/A1 VDD VSS
+ gf180mcu_fd_sc_mcu7t5v0__aoi222_1
XFILLER_61_140 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5831_ hold695/Z _5840_/A2 _5832_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_5762_ _5776_/A1 _5778_/A1 _5762_/A3 _5762_/A4 _5763_/A4 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand4_1
XFILLER_15_590 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_22_538 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_34_387 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4713_ hold85/Z _3819_/Z _4713_/B hold86/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_7501_ _7501_/D _7912_/CLK _7501_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_175_521 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_147_212 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5693_ _5424_/Z _5694_/A4 _5762_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_163_716 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4644_ _4652_/A1 hold61/Z _4644_/B hold62/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_7432_ _7432_/D _7961_/RN _7940_/CLK _7432_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffsnq_1
Xhold712 _7586_/Q hold712/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
X_7363_ _7363_/D _7961_/RN _7565_/CLK _7363_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffsnq_1
X_4575_ hold697/Z _4578_/A2 _4576_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
Xhold701 _7371_/Q hold701/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
X_7294_ _7901_/RN _4334_/Z _7294_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_143_440 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6314_ hold447/Z _6315_/A2 _6315_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
Xhold734 _7878_/Q hold734/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
Xhold745 _7790_/Q hold745/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
Xhold723 _7693_/Q hold723/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
XFILLER_131_613 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_116_676 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xhold767 _7612_/Q hold767/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
Xhold756 _7529_/Q hold756/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
X_6245_ _4448_/Z _6247_/A2 _6245_/B _7756_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_130_134 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_130_123 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_130_112 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6176_ hold675/Z _6191_/A2 _6177_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_5127_ _5648_/A2 _5643_/A2 _5803_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_69_273 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_5058_ _5195_/B _5016_/B _5058_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_85_766 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_29_148 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4009_ _7359_/Q _4488_/A1 _6124_/A1 _7704_/Q _4176_/C _4013_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi221_1
XFILLER_53_652 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_53_641 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_80_460 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_25_354 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_52_162 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_166_510 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_139_702 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_40_368 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_178_392 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_139_757 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_181_524 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_153_215 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_105_2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_4_247 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_136_52 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_134_484 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_122_602 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_96_34 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_453 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
Xhold50 hold50/I hold50/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
XFILLER_76_744 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xhold83 hold83/I hold83/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
Xhold72 hold72/I hold72/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
Xhold61 hold61/I hold61/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
XFILLER_102_392 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xhold94 hold94/I hold94/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
XFILLER_48_479 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_90_235 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_90_224 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_16_321 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_71_471 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_43_184 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XPHY_360 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_176_318 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_31_357 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_129_212 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_84_7 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_61_70 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_8_531 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_177_70 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_8_597 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_8_575 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_99_803 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4360_ _7902_/Q _4360_/A2 _7435_/Q _6623_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_153_771 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_125_484 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_113_602 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_98_302 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_140_421 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4291_ _7973_/Q _4291_/A2 _4291_/B _4292_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi21_2
XFILLER_112_167 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_101_808 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_98_379 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6030_ hold73/Z _6038_/A2 _6030_/B hold183/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_100_318 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_67_744 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
Xclkbuf_0__1040_ _4036_/ZN clkbuf_0__1040_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XTAP_368 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_379 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_20_2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_82_747 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_81_235 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XPHY_19 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_35_641 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6932_ _7914_/Q _7913_/Q _6937_/A1 _6950_/A1 _7195_/C1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor4_4
XFILLER_23_803 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6863_ _7504_/Q _6885_/A2 _6893_/B1 _7389_/Q _6864_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_179_134 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5814_ _4448_/Z _5816_/A2 _5814_/B hold727/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_6794_ _7705_/Q _6889_/A2 _6894_/C1 _7835_/Q _6800_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_148_543 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_5745_ _5579_/B _5804_/A2 _5766_/A2 _5744_/Z _5747_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor4_1
X_5676_ _5747_/A1 _5676_/A2 _5748_/A1 _5676_/B2 _5719_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai22_1
XFILLER_175_373 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4627_ hold79/Z _3830_/Z _4627_/B hold80/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_136_727 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_135_215 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7415_ _7415_/D _7306_/Z _7977_/CLK _7415_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_151_719 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_135_248 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xhold520 _7897_/Q hold520/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
Xhold542 _7459_/Q hold542/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
XFILLER_144_771 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xhold531 _7761_/Q hold531/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
XFILLER_104_602 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_89_302 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
Xhold553 hold553/I _7367_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
X_4558_ _4454_/Z _4558_/A2 _4558_/B _7386_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_7346_ _7346_/D _7301_/Z _7977_/CLK _7346_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
X_7277_ _7277_/A1 _7280_/A2 _7277_/B _7277_/C _7278_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi211_1
Xhold586 hold586/I _7661_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
Xhold597 hold597/I _4783_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
X_4489_ hold762/Z _4504_/A2 _4490_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
Xhold564 _7580_/Q hold564/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
XFILLER_1_228 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
Xhold575 _7400_/Q hold575/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
X_6228_ _4448_/Z _6242_/A2 _6228_/B _7748_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_103_156 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_89_357 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6159_ hold759/Z _6174_/A2 _6160_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_58_744 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_880 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_106_99 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_106_88 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_66_37 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_891 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_18_619 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_72_246 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_122_76 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_72_268 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_53_460 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_81_780 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_13_302 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_41_633 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_53_493 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_158_318 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_13_357 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_182_811 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_31_62 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_181_354 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_31_73 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_31_95 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_147_84 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_147_73 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_135_793 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_110_605 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_49_733 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
Xinput162 wb_sel_i[1] _7281_/C2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
Xinput151 wb_dat_i[30] _7270_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
Xinput140 wb_dat_i[20] _7259_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_163_94 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_76_530 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_49_744 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_76_585 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_64_703 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_36_427 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_64_747 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_17_641 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_63_279 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_51_419 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_44_460 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3860_ _3796_/Z hold133/Z hold134/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_4
XFILLER_16_195 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_20_806 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_177_638 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3791_ _7336_/Q _4383_/A1 _4323_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_31_176 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5530_ _5548_/A2 _5540_/B2 _5530_/B _5803_/A4 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XPHY_190 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
X_5461_ _5461_/A1 _5461_/A2 _5460_/Z _5461_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__and3_1
XFILLER_117_215 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_172_321 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4412_ _7441_/Q input93/Z _7585_/Q _4412_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_68_2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7200_ _7394_/Q _7200_/A2 _7200_/B1 _7388_/Q _7206_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_5392_ _5392_/A1 _5392_/A2 _5376_/B _5405_/B _5392_/B2 _5581_/C VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai32_1
X_4343_ _7520_/Q _4438_/A2 _7515_/Q _4344_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_7131_ _7433_/Q _7936_/Q _7132_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_141_763 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_7062_ _7858_/Q _6938_/I _7188_/A2 _7379_/Q _7063_/A4 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_4274_ _4274_/A1 _4274_/A2 _4274_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_101_638 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_98_176 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6013_ hold73/Z _6021_/A2 _6013_/B hold226/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_79_390 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_39_221 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_39_276 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_36_29 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_7964_ _7964_/D _7317_/Z _7977_/CLK _7964_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XTAP_1309 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_6915_ _6937_/A1 _6953_/A1 _6599_/Z _7197_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor3_4
XFILLER_54_246 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_70_739 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_7895_ _7895_/D _7901_/RN _7895_/CLK _7895_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_63_780 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_23_611 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_168_605 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6846_ _7755_/Q _6644_/Z _6885_/B1 _7715_/Q _6847_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_167_115 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6777_ _6777_/A1 _6777_/A2 _6777_/A3 _6778_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor3_1
XFILLER_22_176 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_50_463 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5728_ _5287_/C _5316_/B _5762_/A4 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_3989_ _3989_/A1 _3989_/A2 _3989_/A3 _3989_/A4 _3990_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand4_2
XFILLER_22_187 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_182_107 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_176_671 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5659_ _5674_/A1 _5674_/A2 _5657_/Z _5674_/A3 _5675_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand4_1
XFILLER_163_354 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_117_771 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_2_515 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_144_590 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_132_741 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_117_793 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
Xhold361 _7857_/Q hold361/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
XFILLER_89_121 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
Xhold350 _7449_/Q hold350/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
X_7329_ input75/Z _4334_/Z _7329_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__and2_1
Xhold394 hold394/I _7674_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
Xhold383 hold383/I _7658_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
Xhold372 _7881_/Q hold372/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
XFILLER_89_198 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_92_308 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_18_416 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_46_703 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_172_2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_133_86 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_100_682 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_73_522 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_46_747 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_93_79 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_73_566 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1843 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1832 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1821 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1810 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_26_460 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1876 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1865 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1854 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_159_649 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_159_638 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1898 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1887 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_41_463 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_154_321 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_182_674 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_123_763 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_150_593 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_123_785 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_1_570 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_3_88 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_91_363 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4961_ _5022_/B _4944_/Z _4963_/A4 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_64_588 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_45_780 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3912_ _7691_/Q _6090_/A1 _6158_/A1 _7723_/Q _3916_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_7680_ _7680_/D _7961_/RN _7815_/CLK _7680_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
X_6700_ _7717_/Q _6881_/A2 _6882_/B1 _7653_/Q _6702_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_4892_ _4454_/Z _4892_/A2 _4892_/B _7536_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_3843_ _3801_/Z _3864_/A2 _3843_/A3 hold274/Z _4075_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand4_4
X_6631_ _7909_/Q _7908_/Q _6662_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_4
XFILLER_32_463 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_177_479 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_158_660 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_118_513 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6562_ _6562_/A1 _6561_/Z _6564_/B _6563_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_3774_ _7345_/Q _3774_/A2 _3763_/B _3774_/B _7965_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai31_1
XFILLER_173_641 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_5513_ _5179_/B _5793_/A2 _5555_/B _5514_/A4 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_6493_ hold529/Z _6502_/A2 _6494_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_161_803 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_145_354 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5444_ _5627_/A2 _5444_/A2 _5613_/A2 _5444_/A4 _5445_/A4 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand4_1
X_5375_ _5015_/B _5197_/Z _5375_/A3 _5375_/A4 _5708_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor4_4
XFILLER_99_463 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7114_ _7900_/Q _7197_/A2 _7196_/A2 _7892_/Q _7196_/B1 _7642_/Q _7116_/A3 VDD VSS
+ gf180mcu_fd_sc_mcu7t5v0__aoi222_1
XFILLER_101_424 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_59_327 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4326_ _7411_/Q _3738_/Z _4327_/S VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_7045_ _7761_/Q _7202_/C2 _7205_/A2 _7735_/Q _7048_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_4257_ _7504_/Q _4831_/A1 hold21/I _4215_/Z _4260_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_170_29 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_86_179 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4188_ _7863_/Q _6469_/A1 _4554_/A1 _7386_/Q _7356_/Q _4488_/A1 _4203_/A2 VDD VSS
+ gf180mcu_fd_sc_mcu7t5v0__aoi222_2
XFILLER_67_371 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_28_747 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_55_511 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_103_89 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_82_396 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7947_ _7947_/D _7949_/CLK _7947_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_70_514 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1117 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1128 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1106 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_43_739 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_7878_ _7878_/D _7901_/RN _7890_/CLK _7878_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffsnq_1
XTAP_1139 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_6829_ _7133_/S _6829_/A2 _6829_/B _7927_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_51_783 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_168_479 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_10_124 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_23_496 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_23_485 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_149_682 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_148_170 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_136_321 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_10_179 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_164_685 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_88_46 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_151_357 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xhold180 hold180/I _7856_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
XFILLER_2_334 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xhold191 _7747_/Q hold191/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
XFILLER_132_582 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_105_785 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_2_389 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_120_755 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_144_96 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_92_105 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_77_168 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_19_703 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_92_149 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_86_680 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_19_747 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2352 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2341 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2330 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2396 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2385 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2374 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2363 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1651 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1640 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1684 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1673 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1662 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_14_463 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1695 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_41_282 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_169_93 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_155_641 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_143_803 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_127_354 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_115_549 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5160_ _5538_/A1 _5390_/A2 _5162_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_123_582 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5091_ _5058_/Z _5456_/A2 _5114_/A3 _5579_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__and3_2
XFILLER_110_210 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4111_ _3817_/I hold25/Z _5881_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_2
XFILLER_110_254 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4042_ _7793_/Q _6316_/A1 _4067_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_84_617 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_84_628 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_68_179 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_83_138 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_7801_ _7801_/D _7901_/RN _7868_/CLK _7801_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_80_812 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_64_374 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_5993_ hold175/Z _6004_/A2 hold176/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_178_700 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4944_ _5338_/A1 _4900_/Z _4944_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__xor2_2
XFILLER_40_709 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7732_ _7732_/D _7961_/RN _7733_/CLK _7732_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffsnq_1
XFILLER_178_744 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_33_783 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7663_ _7663_/D _7901_/RN _7812_/CLK _7663_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
X_4875_ _4448_/Z _4877_/A2 _4875_/B _7529_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_7594_ _7594_/D _7901_/RN _7865_/CLK _8004_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
X_3826_ hold124/Z _4153_/A1 _5954_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_4
X_6614_ _6953_/A2 _6950_/A2 _6955_/A4 _7193_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor3_4
XFILLER_118_321 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_6545_ hold73/Z _6553_/A2 _6545_/B _7897_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_3757_ _3765_/A1 _3765_/A2 _3762_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_161_611 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3688_ _7793_/Q _3688_/ZN VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_106_538 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6476_ hold364/Z _6485_/A2 _6477_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
Xoutput230 _8003_/Z mgmt_gpio_out[29] VDD VSS gf180mcu_fd_sc_mcu7t5v0__buf_8
XFILLER_133_357 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5427_ _5685_/B _5247_/B _5540_/C _5686_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi21_1
Xoutput252 _4422_/ZN pad_flash_io0_ie VDD VSS gf180mcu_fd_sc_mcu7t5v0__buf_8
Xoutput241 _7985_/Z mgmt_gpio_out[4] VDD VSS gf180mcu_fd_sc_mcu7t5v0__buf_8
XFILLER_160_187 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_160_176 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5358_ _5741_/A1 _5602_/A1 _5741_/A3 _5636_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor3_2
XFILLER_102_700 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
Xoutput263 _7559_/Q pll_div[1] VDD VSS gf180mcu_fd_sc_mcu7t5v0__buf_8
Xoutput274 _7359_/Q pll_trim[12] VDD VSS gf180mcu_fd_sc_mcu7t5v0__buf_8
Xoutput285 _7353_/Q pll_trim[22] VDD VSS gf180mcu_fd_sc_mcu7t5v0__buf_8
X_4309_ _4308_/Z _7340_/Q _4309_/S _7340_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_102_744 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_59_124 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
Xoutput296 _7356_/Q pll_trim[9] VDD VSS gf180mcu_fd_sc_mcu7t5v0__buf_8
X_5289_ _3723_/I _5579_/B _5721_/C _5680_/C _5293_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XFILLER_114_33 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7028_ _7433_/Q _7932_/Q _7028_/B _7030_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_59_157 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_114_44 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_102_799 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_87_499 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_83_661 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_74_37 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_71_812 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_43_503 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_43_514 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_168_210 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_90_25 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_23_282 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_135_2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_137_641 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_11_499 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_11_488 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_164_460 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_109_354 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_99_56 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_99_34 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_124_313 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_99_67 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_155_73 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_97_208 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_3_698 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_709 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_155_95 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_151_198 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_93_425 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_93_458 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_81_609 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_34 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_46_330 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_80_108 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_62_812 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2171 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2160 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_46_396 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
Xnet299_2 net299_2/I _4416_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XTAP_2193 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2182 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_21_219 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1492 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1481 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1470 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_14_271 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_15_783 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_30_720 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_175_736 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4660_ _7459_/Q hold55/I hold36/Z hold37/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_9_98 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6330_ hold68/Z _6332_/A2 _6330_/B hold288/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_128_663 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_4591_ _4448_/Z _4593_/A2 _4591_/B _7399_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_143_611 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_127_184 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_50_2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6261_ hold460/Z _6264_/A2 _6262_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_115_357 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_89_709 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5212_ _4906_/Z _5373_/A3 _5373_/A4 _5212_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__and3_1
XFILLER_170_463 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6192_ _6192_/A1 hold32/Z _6208_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_4
XFILLER_103_519 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8000_ _8000_/I _8000_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_5143_ _5645_/A1 _5545_/A2 _5768_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_142_187 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_5074_ _5600_/A1 _5797_/B _5783_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_4
XFILLER_69_499 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_56_105 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_56_138 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4025_ _4025_/A1 _4025_/A2 _4025_/A3 _4025_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__or3_1
XFILLER_44_29 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5976_ hold249/Z _5987_/A2 _5977_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_13_709 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4927_ _5211_/A3 _4920_/Z _5011_/B _4951_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi21_2
X_7715_ _7715_/D _7901_/RN _7812_/CLK _7715_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_100_24 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_33_580 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_166_703 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7646_ hold30/Z _7961_/RN _7706_/CLK _7646_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffsnq_1
X_4858_ _4858_/A1 _7285_/A2 _4862_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_178_596 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_166_747 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3809_ _7506_/Q hold23/Z _3811_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_121_8 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_181_728 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_119_641 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_109_22 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4789_ _7480_/Q _4795_/S _4790_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_7577_ _7577_/D _7961_/RN _7645_/CLK _7577_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_146_460 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6528_ hold73/Z _6536_/A2 _6528_/B _7889_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_109_66 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6459_ hold361/Z _6468_/A2 _6460_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
Xclkbuf_leaf_7_csclk clkbuf_leaf_9_csclk/I _7834_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_133_176 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_624 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_75_436 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_75_458 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_18_41 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_62_108 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_28_363 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_44_812 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_55_160 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_16_558 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_43_344 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_169_552 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_24_580 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_11_241 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_157_769 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_7_212 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_144_419 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_165_780 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_166_72 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_152_463 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_112_305 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_112_316 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_506 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_112_327 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_79_753 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_539 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_528 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_517 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_38_105 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_66_458 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_81_428 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_35_812 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_47_672 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_62_620 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5830_ _4448_/Z _5840_/A2 _5830_/B _7563_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_22_517 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5761_ _5686_/Z _5761_/A2 _5758_/Z _5760_/Z _5786_/B1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand4_1
XFILLER_98_2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_61_174 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4712_ _3819_/Z hold68/Z _4713_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_7500_ _7500_/D _7949_/CLK _7500_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_5692_ _5692_/A1 _5692_/A2 _5692_/B _5694_/A4 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_148_747 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7431_ hold99/Z _7901_/RN _7603_/CLK hold97/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_175_566 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4643_ hold60/Z _3830_/Z _4643_/B hold61/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_135_419 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_128_460 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_116_600 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
Xhold702 _7364_/Q hold702/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
X_7362_ _7362_/D _7961_/RN _7875_/CLK _7362_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffsnq_2
X_4574_ _4574_/A1 _7285_/A2 _4578_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_7293_ _7901_/RN _4334_/Z _7293_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_116_633 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6313_ hold68/Z _6315_/A2 _6313_/B _7788_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
Xhold713 _7685_/Q hold713/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
Xhold735 _7348_/Q hold735/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
Xhold746 _7636_/Q hold746/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
Xhold724 _7444_/Q hold724/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
XFILLER_171_783 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
Xhold768 _7652_/Q hold768/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
Xhold757 _7960_/Q hold757/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
X_6244_ hold654/Z _6247_/A2 _6245_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_170_282 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_143_496 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_39_29 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_6175_ hold119/Z hold32/Z _6191_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_4
XFILLER_85_712 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_85_701 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_5126_ _5390_/A2 _5122_/Z _5479_/A2 _5669_/A1 _5651_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_130_179 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_69_263 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_29_105 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_57_425 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5057_ _5303_/A3 _5421_/A1 _5319_/C VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_4
XFILLER_85_778 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_84_277 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4008_ _7624_/Q _5954_/A1 _4020_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_26_812 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_38_672 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_44_108 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_65_491 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_25_366 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_52_130 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_5959_ hold184/Z _5970_/A2 hold185/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_40_325 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_52_174 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_53_697 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_154_717 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_7629_ _7629_/D _7901_/RN _7797_/CLK _7629_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffsnq_1
XFILLER_138_257 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_181_514 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_153_227 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_153_205 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_147_780 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_4_204 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_106_132 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_134_463 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_121_102 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_106_176 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_96_46 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
Xhold40 hold40/I hold40/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
Xhold73 hold73/I hold73/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
Xhold62 hold62/I hold62/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
Xhold51 hold51/I hold51/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
XFILLER_29_73 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xhold95 hold95/I hold95/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
Xhold84 hold84/I hold84/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
XFILLER_63_428 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_17_812 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_91_759 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_90_247 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_56_480 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_56_491 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_90_269 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_90_258 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_43_141 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_43_130 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_45_50 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XPHY_361 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_350 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_145_706 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_61_82 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_145_739 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_6_44 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_153_783 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_140_400 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_125_496 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4290_ _7973_/Q _4291_/A2 _4382_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_112_157 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_112_179 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_67_712 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_369 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_39_425 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_94_553 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_94_531 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_66_233 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_13_2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_26_108 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_7980_ _7980_/D _7333_/Z _4418_/I1 _7980_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_81_247 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6931_ _6937_/A1 _6941_/A1 _7196_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_4
X_6862_ _7405_/Q _6883_/A2 _6883_/B1 _7397_/Q _6864_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_168_809 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5813_ hold726/Z _5816_/A2 _5814_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_6793_ _7641_/Q _6890_/A2 _6665_/Z _7745_/Q _6793_/C _6800_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi221_1
XFILLER_148_522 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_5744_ _5499_/Z _5542_/Z _5744_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__or2_1
XFILLER_148_555 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5675_ _5675_/A1 _5671_/Z _5676_/B2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_1
Xclkbuf_leaf_72_csclk _7961_/CLK _7960_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
X_4626_ _3830_/Z _4454_/Z _4627_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_135_205 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_7414_ _7414_/D _7305_/Z _4418_/I1 _7414_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_4
XFILLER_151_709 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_135_238 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
Xhold510 _7788_/Q hold510/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
X_7345_ _7345_/D _7300_/Z _7977_/CLK _7345_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_2
XFILLER_116_463 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xhold521 _7787_/Q hold521/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
Xhold532 _7369_/Q hold532/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
Xhold543 _7368_/Q hold543/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
Xhold554 _7567_/Q hold554/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
X_4557_ hold632/Z _4558_/A2 _4558_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_7276_ _7276_/A1 _7276_/A2 _7277_/C VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
Xhold565 _7709_/Q hold565/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
XFILLER_104_636 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
Xhold587 _7495_/Q hold587/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
X_4488_ _4488_/A1 _7285_/A2 _4504_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_4
Xclkbuf_leaf_87_csclk _7396_/CLK _7572_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
Xhold576 _7408_/Q hold576/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
X_6227_ hold650/Z _6242_/A2 _6228_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_131_444 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_106_34 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_58_701 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xhold598 hold598/I _7477_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
XFILLER_131_499 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6158_ _6158_/A1 hold32/Z _6174_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_4
XTAP_870 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_5109_ _5669_/A1 _5672_/A2 _5673_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
Xclkbuf_leaf_10_csclk clkbuf_leaf_9_csclk/I _7826_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XTAP_881 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_892 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_6089_ hold90/Z _6089_/A2 _6089_/B hold239/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_57_266 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_122_33 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_38_480 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_45_428 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_57_288 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xclkbuf_leaf_25_csclk _7825_/CLK _7868_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_82_37 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_25_141 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_159_809 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_81_770 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_26_697 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_21_380 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_127_739 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_181_366 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_135_783 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_135_772 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_150_742 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_134_282 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_107_496 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_150_764 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_163_73 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_163_62 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_251 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_1_785 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_49_712 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xinput163 wb_sel_i[2] _7281_/B1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
Xinput152 wb_dat_i[31] _7275_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
Xinput141 wb_dat_i[21] _7265_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
Xinput130 wb_dat_i[11] _7255_/B1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_163_84 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_49_789 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_91_567 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_44_450 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_176_105 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_176_127 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_3790_ hold126/Z _3789_/Z _3810_/S _3790_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_4
XFILLER_72_92 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_31_144 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_191 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_180 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
X_5460_ _5460_/A1 _5460_/A2 _5657_/A3 _5460_/A4 _5460_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__and4_1
X_4411_ _7442_/Q _4411_/I1 _7583_/Q _4411_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_133_709 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_126_761 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_99_601 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5391_ _5741_/A1 _4993_/B _5797_/A1 _5391_/B _5735_/C VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai31_1
X_4342_ _4342_/I _7519_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_113_400 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7130_ _7130_/A1 _7130_/A2 _7130_/A3 _6949_/I _7610_/Q _7132_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai32_1
XFILLER_98_155 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7061_ _7648_/Q _7195_/A2 _7195_/B1 _7624_/Q _7195_/C1 _7874_/Q _7063_/A3 VDD VSS
+ gf180mcu_fd_sc_mcu7t5v0__aoi222_1
X_4273_ _7563_/Q _5828_/A1 _4574_/A1 _7393_/Q _4274_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_141_797 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_140_263 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_113_499 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_113_488 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_98_166 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_6012_ hold224/Z _6021_/A2 hold225/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
.ends

