VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO mprj_io_buffer
  CLASS BLOCK ;
  FOREIGN mprj_io_buffer ;
  ORIGIN 0.000 0.000 ;
  SIZE 85.000 BY 60.000 ;
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER Metal4 ;
        RECT 10.610 7.540 12.210 51.260 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 31.190 7.540 32.790 51.260 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 51.770 7.540 53.370 51.260 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 72.350 7.540 73.950 51.260 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER Metal4 ;
        RECT 20.900 7.540 22.500 51.260 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 41.480 7.540 43.080 51.260 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 62.060 7.540 63.660 51.260 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 82.640 7.540 84.240 51.260 ;
    END
  END VSS
  PIN mgmt_gpio_in[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 2.800 0.000 3.360 4.000 ;
    END
  END mgmt_gpio_in[0]
  PIN mgmt_gpio_in[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 25.200 0.000 25.760 4.000 ;
    END
  END mgmt_gpio_in[10]
  PIN mgmt_gpio_in[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 27.440 0.000 28.000 4.000 ;
    END
  END mgmt_gpio_in[11]
  PIN mgmt_gpio_in[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 29.680 0.000 30.240 4.000 ;
    END
  END mgmt_gpio_in[12]
  PIN mgmt_gpio_in[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 31.920 0.000 32.480 4.000 ;
    END
  END mgmt_gpio_in[13]
  PIN mgmt_gpio_in[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 34.160 0.000 34.720 4.000 ;
    END
  END mgmt_gpio_in[14]
  PIN mgmt_gpio_in[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 36.400 0.000 36.960 4.000 ;
    END
  END mgmt_gpio_in[15]
  PIN mgmt_gpio_in[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 38.640 0.000 39.200 4.000 ;
    END
  END mgmt_gpio_in[16]
  PIN mgmt_gpio_in[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 40.880 0.000 41.440 4.000 ;
    END
  END mgmt_gpio_in[17]
  PIN mgmt_gpio_in[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 5.040 0.000 5.600 4.000 ;
    END
  END mgmt_gpio_in[1]
  PIN mgmt_gpio_in[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 7.280 0.000 7.840 4.000 ;
    END
  END mgmt_gpio_in[2]
  PIN mgmt_gpio_in[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 9.520 0.000 10.080 4.000 ;
    END
  END mgmt_gpio_in[3]
  PIN mgmt_gpio_in[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 11.760 0.000 12.320 4.000 ;
    END
  END mgmt_gpio_in[4]
  PIN mgmt_gpio_in[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 14.000 0.000 14.560 4.000 ;
    END
  END mgmt_gpio_in[5]
  PIN mgmt_gpio_in[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 16.240 0.000 16.800 4.000 ;
    END
  END mgmt_gpio_in[6]
  PIN mgmt_gpio_in[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 18.480 0.000 19.040 4.000 ;
    END
  END mgmt_gpio_in[7]
  PIN mgmt_gpio_in[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 20.720 0.000 21.280 4.000 ;
    END
  END mgmt_gpio_in[8]
  PIN mgmt_gpio_in[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 22.960 0.000 23.520 4.000 ;
    END
  END mgmt_gpio_in[9]
  PIN mgmt_gpio_in_buf[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 2.800 56.000 3.360 60.000 ;
    END
  END mgmt_gpio_in_buf[0]
  PIN mgmt_gpio_in_buf[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 25.200 56.000 25.760 60.000 ;
    END
  END mgmt_gpio_in_buf[10]
  PIN mgmt_gpio_in_buf[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 27.440 56.000 28.000 60.000 ;
    END
  END mgmt_gpio_in_buf[11]
  PIN mgmt_gpio_in_buf[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 29.680 56.000 30.240 60.000 ;
    END
  END mgmt_gpio_in_buf[12]
  PIN mgmt_gpio_in_buf[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 31.920 56.000 32.480 60.000 ;
    END
  END mgmt_gpio_in_buf[13]
  PIN mgmt_gpio_in_buf[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 34.160 56.000 34.720 60.000 ;
    END
  END mgmt_gpio_in_buf[14]
  PIN mgmt_gpio_in_buf[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 36.400 56.000 36.960 60.000 ;
    END
  END mgmt_gpio_in_buf[15]
  PIN mgmt_gpio_in_buf[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 38.640 56.000 39.200 60.000 ;
    END
  END mgmt_gpio_in_buf[16]
  PIN mgmt_gpio_in_buf[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 40.880 56.000 41.440 60.000 ;
    END
  END mgmt_gpio_in_buf[17]
  PIN mgmt_gpio_in_buf[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 5.040 56.000 5.600 60.000 ;
    END
  END mgmt_gpio_in_buf[1]
  PIN mgmt_gpio_in_buf[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 7.280 56.000 7.840 60.000 ;
    END
  END mgmt_gpio_in_buf[2]
  PIN mgmt_gpio_in_buf[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 9.520 56.000 10.080 60.000 ;
    END
  END mgmt_gpio_in_buf[3]
  PIN mgmt_gpio_in_buf[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 11.760 56.000 12.320 60.000 ;
    END
  END mgmt_gpio_in_buf[4]
  PIN mgmt_gpio_in_buf[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 14.000 56.000 14.560 60.000 ;
    END
  END mgmt_gpio_in_buf[5]
  PIN mgmt_gpio_in_buf[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 16.240 56.000 16.800 60.000 ;
    END
  END mgmt_gpio_in_buf[6]
  PIN mgmt_gpio_in_buf[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 18.480 56.000 19.040 60.000 ;
    END
  END mgmt_gpio_in_buf[7]
  PIN mgmt_gpio_in_buf[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 20.720 56.000 21.280 60.000 ;
    END
  END mgmt_gpio_in_buf[8]
  PIN mgmt_gpio_in_buf[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 22.960 56.000 23.520 60.000 ;
    END
  END mgmt_gpio_in_buf[9]
  PIN mgmt_gpio_oeb[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 14.560 4.000 15.120 ;
    END
  END mgmt_gpio_oeb[0]
  PIN mgmt_gpio_oeb[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 44.240 4.000 44.800 ;
    END
  END mgmt_gpio_oeb[1]
  PIN mgmt_gpio_oeb_buf[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 81.000 14.560 85.000 15.120 ;
    END
  END mgmt_gpio_oeb_buf[0]
  PIN mgmt_gpio_oeb_buf[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 81.000 44.240 85.000 44.800 ;
    END
  END mgmt_gpio_oeb_buf[1]
  PIN mgmt_gpio_out[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 43.120 56.000 43.680 60.000 ;
    END
  END mgmt_gpio_out[0]
  PIN mgmt_gpio_out[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 65.520 56.000 66.080 60.000 ;
    END
  END mgmt_gpio_out[10]
  PIN mgmt_gpio_out[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 67.760 56.000 68.320 60.000 ;
    END
  END mgmt_gpio_out[11]
  PIN mgmt_gpio_out[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 70.000 56.000 70.560 60.000 ;
    END
  END mgmt_gpio_out[12]
  PIN mgmt_gpio_out[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 72.240 56.000 72.800 60.000 ;
    END
  END mgmt_gpio_out[13]
  PIN mgmt_gpio_out[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 74.480 56.000 75.040 60.000 ;
    END
  END mgmt_gpio_out[14]
  PIN mgmt_gpio_out[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 76.720 56.000 77.280 60.000 ;
    END
  END mgmt_gpio_out[15]
  PIN mgmt_gpio_out[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 78.960 56.000 79.520 60.000 ;
    END
  END mgmt_gpio_out[16]
  PIN mgmt_gpio_out[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 81.200 56.000 81.760 60.000 ;
    END
  END mgmt_gpio_out[17]
  PIN mgmt_gpio_out[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 45.360 56.000 45.920 60.000 ;
    END
  END mgmt_gpio_out[1]
  PIN mgmt_gpio_out[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 47.600 56.000 48.160 60.000 ;
    END
  END mgmt_gpio_out[2]
  PIN mgmt_gpio_out[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 49.840 56.000 50.400 60.000 ;
    END
  END mgmt_gpio_out[3]
  PIN mgmt_gpio_out[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 52.080 56.000 52.640 60.000 ;
    END
  END mgmt_gpio_out[4]
  PIN mgmt_gpio_out[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 54.320 56.000 54.880 60.000 ;
    END
  END mgmt_gpio_out[5]
  PIN mgmt_gpio_out[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 56.560 56.000 57.120 60.000 ;
    END
  END mgmt_gpio_out[6]
  PIN mgmt_gpio_out[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 58.800 56.000 59.360 60.000 ;
    END
  END mgmt_gpio_out[7]
  PIN mgmt_gpio_out[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 61.040 56.000 61.600 60.000 ;
    END
  END mgmt_gpio_out[8]
  PIN mgmt_gpio_out[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 63.280 56.000 63.840 60.000 ;
    END
  END mgmt_gpio_out[9]
  PIN mgmt_gpio_out_buf[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 43.120 0.000 43.680 4.000 ;
    END
  END mgmt_gpio_out_buf[0]
  PIN mgmt_gpio_out_buf[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 65.520 0.000 66.080 4.000 ;
    END
  END mgmt_gpio_out_buf[10]
  PIN mgmt_gpio_out_buf[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 67.760 0.000 68.320 4.000 ;
    END
  END mgmt_gpio_out_buf[11]
  PIN mgmt_gpio_out_buf[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 70.000 0.000 70.560 4.000 ;
    END
  END mgmt_gpio_out_buf[12]
  PIN mgmt_gpio_out_buf[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 72.240 0.000 72.800 4.000 ;
    END
  END mgmt_gpio_out_buf[13]
  PIN mgmt_gpio_out_buf[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 74.480 0.000 75.040 4.000 ;
    END
  END mgmt_gpio_out_buf[14]
  PIN mgmt_gpio_out_buf[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 76.720 0.000 77.280 4.000 ;
    END
  END mgmt_gpio_out_buf[15]
  PIN mgmt_gpio_out_buf[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 78.960 0.000 79.520 4.000 ;
    END
  END mgmt_gpio_out_buf[16]
  PIN mgmt_gpio_out_buf[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 81.200 0.000 81.760 4.000 ;
    END
  END mgmt_gpio_out_buf[17]
  PIN mgmt_gpio_out_buf[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 45.360 0.000 45.920 4.000 ;
    END
  END mgmt_gpio_out_buf[1]
  PIN mgmt_gpio_out_buf[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 47.600 0.000 48.160 4.000 ;
    END
  END mgmt_gpio_out_buf[2]
  PIN mgmt_gpio_out_buf[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 49.840 0.000 50.400 4.000 ;
    END
  END mgmt_gpio_out_buf[3]
  PIN mgmt_gpio_out_buf[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 52.080 0.000 52.640 4.000 ;
    END
  END mgmt_gpio_out_buf[4]
  PIN mgmt_gpio_out_buf[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 54.320 0.000 54.880 4.000 ;
    END
  END mgmt_gpio_out_buf[5]
  PIN mgmt_gpio_out_buf[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 56.560 0.000 57.120 4.000 ;
    END
  END mgmt_gpio_out_buf[6]
  PIN mgmt_gpio_out_buf[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 58.800 0.000 59.360 4.000 ;
    END
  END mgmt_gpio_out_buf[7]
  PIN mgmt_gpio_out_buf[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 61.040 0.000 61.600 4.000 ;
    END
  END mgmt_gpio_out_buf[8]
  PIN mgmt_gpio_out_buf[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 63.280 0.000 63.840 4.000 ;
    END
  END mgmt_gpio_out_buf[9]
  OBS
      LAYER Metal1 ;
        RECT 1.120 7.540 84.240 51.260 ;
      LAYER Metal2 ;
        RECT 3.660 55.700 4.740 56.000 ;
        RECT 5.900 55.700 6.980 56.000 ;
        RECT 8.140 55.700 9.220 56.000 ;
        RECT 10.380 55.700 11.460 56.000 ;
        RECT 12.620 55.700 13.700 56.000 ;
        RECT 14.860 55.700 15.940 56.000 ;
        RECT 17.100 55.700 18.180 56.000 ;
        RECT 19.340 55.700 20.420 56.000 ;
        RECT 21.580 55.700 22.660 56.000 ;
        RECT 23.820 55.700 24.900 56.000 ;
        RECT 26.060 55.700 27.140 56.000 ;
        RECT 28.300 55.700 29.380 56.000 ;
        RECT 30.540 55.700 31.620 56.000 ;
        RECT 32.780 55.700 33.860 56.000 ;
        RECT 35.020 55.700 36.100 56.000 ;
        RECT 37.260 55.700 38.340 56.000 ;
        RECT 39.500 55.700 40.580 56.000 ;
        RECT 41.740 55.700 42.820 56.000 ;
        RECT 43.980 55.700 45.060 56.000 ;
        RECT 46.220 55.700 47.300 56.000 ;
        RECT 48.460 55.700 49.540 56.000 ;
        RECT 50.700 55.700 51.780 56.000 ;
        RECT 52.940 55.700 54.020 56.000 ;
        RECT 55.180 55.700 56.260 56.000 ;
        RECT 57.420 55.700 58.500 56.000 ;
        RECT 59.660 55.700 60.740 56.000 ;
        RECT 61.900 55.700 62.980 56.000 ;
        RECT 64.140 55.700 65.220 56.000 ;
        RECT 66.380 55.700 67.460 56.000 ;
        RECT 68.620 55.700 69.700 56.000 ;
        RECT 70.860 55.700 71.940 56.000 ;
        RECT 73.100 55.700 74.180 56.000 ;
        RECT 75.340 55.700 76.420 56.000 ;
        RECT 77.580 55.700 78.660 56.000 ;
        RECT 79.820 55.700 80.900 56.000 ;
        RECT 82.060 55.700 84.100 56.000 ;
        RECT 2.940 4.300 84.100 55.700 ;
        RECT 3.660 4.000 4.740 4.300 ;
        RECT 5.900 4.000 6.980 4.300 ;
        RECT 8.140 4.000 9.220 4.300 ;
        RECT 10.380 4.000 11.460 4.300 ;
        RECT 12.620 4.000 13.700 4.300 ;
        RECT 14.860 4.000 15.940 4.300 ;
        RECT 17.100 4.000 18.180 4.300 ;
        RECT 19.340 4.000 20.420 4.300 ;
        RECT 21.580 4.000 22.660 4.300 ;
        RECT 23.820 4.000 24.900 4.300 ;
        RECT 26.060 4.000 27.140 4.300 ;
        RECT 28.300 4.000 29.380 4.300 ;
        RECT 30.540 4.000 31.620 4.300 ;
        RECT 32.780 4.000 33.860 4.300 ;
        RECT 35.020 4.000 36.100 4.300 ;
        RECT 37.260 4.000 38.340 4.300 ;
        RECT 39.500 4.000 40.580 4.300 ;
        RECT 41.740 4.000 42.820 4.300 ;
        RECT 43.980 4.000 45.060 4.300 ;
        RECT 46.220 4.000 47.300 4.300 ;
        RECT 48.460 4.000 49.540 4.300 ;
        RECT 50.700 4.000 51.780 4.300 ;
        RECT 52.940 4.000 54.020 4.300 ;
        RECT 55.180 4.000 56.260 4.300 ;
        RECT 57.420 4.000 58.500 4.300 ;
        RECT 59.660 4.000 60.740 4.300 ;
        RECT 61.900 4.000 62.980 4.300 ;
        RECT 64.140 4.000 65.220 4.300 ;
        RECT 66.380 4.000 67.460 4.300 ;
        RECT 68.620 4.000 69.700 4.300 ;
        RECT 70.860 4.000 71.940 4.300 ;
        RECT 73.100 4.000 74.180 4.300 ;
        RECT 75.340 4.000 76.420 4.300 ;
        RECT 77.580 4.000 78.660 4.300 ;
        RECT 79.820 4.000 80.900 4.300 ;
        RECT 82.060 4.000 84.100 4.300 ;
      LAYER Metal3 ;
        RECT 2.890 45.100 84.150 51.100 ;
        RECT 4.300 43.940 80.700 45.100 ;
        RECT 2.890 15.420 84.150 43.940 ;
        RECT 4.300 14.260 80.700 15.420 ;
        RECT 2.890 7.700 84.150 14.260 ;
  END
END mprj_io_buffer
END LIBRARY

