* NGSPICE file created from housekeeping.ext - technology: gf180mcuC

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__fill_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__fill_2 VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__fillcap_4 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__fillcap_4 VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__dffnsnq_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__dffnsnq_1 D SETN CLKN Q VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__fill_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__fill_1 VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__nor2_4 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__nor2_4 A1 A2 ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__dffsnq_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__dffsnq_1 D SETN CLK Q VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__aoi222_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__aoi222_1 A1 A2 B1 B2 C1 C2 ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__aoi22_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__aoi22_1 A1 A2 B1 B2 ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__nand4_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__nand4_1 A1 A2 A3 A4 ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__nand4_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__nand4_2 A1 A2 A3 A4 ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__fillcap_8 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__fillcap_8 VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__oai21_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__oai21_1 A1 A2 B ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__nor3_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__nor3_1 A1 A2 A3 ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__nand2_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__nand2_1 A1 A2 ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__and2_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__and2_1 A1 A2 Z VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__dlyd_4 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__dlyd_4 I Z VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__fillcap_16 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__fillcap_16 VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__filltie abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__filltie VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__or2_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__or2_1 A1 A2 Z VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__nand2_4 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__nand2_4 A1 A2 ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__aoi21_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__aoi21_1 A1 A2 B ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__aoi211_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__aoi211_1 A1 A2 B C ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__nor2_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__nor2_1 A1 A2 ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__nor4_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__nor4_2 A1 A2 A3 A4 ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__dffq_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__dffq_1 D CLK Q VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 D RN CLK Q VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__nor2_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__nor2_2 A1 A2 ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__mux2_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__mux2_2 I0 I1 S Z VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__xor2_4 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__xor2_4 A1 A2 Z VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__oai31_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__oai31_2 A1 A2 A3 B ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__clkinv_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__clkinv_1 I ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__buf_4 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__buf_4 I Z VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__nand4_4 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__nand4_4 A1 A2 A3 A4 ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__or4_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__or4_2 A1 A2 A3 A4 Z VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__oai22_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__oai22_1 A1 A2 B1 B2 ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__and3_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__and3_1 A1 A2 A3 Z VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__nor4_4 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__nor4_4 A1 A2 A3 A4 ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 I Z VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__endcap abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__endcap VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__fillcap_32 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__fillcap_32 VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__nand3_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__nand3_1 A1 A2 A3 ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__dffrnq_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__dffrnq_2 D RN CLK Q VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__nor3_4 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__nor3_4 A1 A2 A3 ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__buf_12 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__buf_12 I Z VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__dlyb_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__dlyb_1 I Z VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__dffnrnq_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__dffnrnq_1 D RN CLKN Q VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__nand3_4 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__nand3_4 A1 A2 A3 ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__and4_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__and4_1 A1 A2 A3 A4 Z VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__aoi221_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__aoi221_1 A1 A2 B1 B2 C ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__oai32_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__oai32_1 A1 A2 A3 B1 B2 ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__oai21_4 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__oai21_4 A1 A2 B ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__oai21_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__oai21_2 A1 A2 B ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__nor4_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__nor4_1 A1 A2 A3 A4 ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__oai211_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__oai211_1 A1 A2 B C ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__or2_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__or2_2 A1 A2 Z VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__nand2_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__nand2_2 A1 A2 ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__nor3_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__nor3_2 A1 A2 A3 ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__buf_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__buf_2 I Z VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__aoi211_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__aoi211_2 A1 A2 B C ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__aoi211_4 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__aoi211_4 A1 A2 B C ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__xor2_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__xor2_1 A1 A2 Z VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__aoi21_4 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__aoi21_4 A1 A2 B ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__oai31_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__oai31_1 A1 A2 A3 B ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__dffsnq_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__dffsnq_2 D SETN CLK Q VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__dlyc_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__dlyc_1 I Z VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__buf_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__buf_1 I Z VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__dffrnq_4 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__dffrnq_4 D RN CLK Q VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__or3_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__or3_1 A1 A2 A3 Z VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__clkinv_3 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__clkinv_3 I ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__or4_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__or4_1 A1 A2 A3 A4 Z VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__dlyd_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__dlyd_1 I Z VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__inv_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__inv_2 I ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__clkbuf_12 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__clkbuf_12 I Z VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__aoi222_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__aoi222_2 A1 A2 B1 B2 C1 C2 ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__or2_4 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__or2_4 A1 A2 Z VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__or3_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__or3_2 A1 A2 A3 Z VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__dffsnq_4 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__dffsnq_4 D SETN CLK Q VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__clkinv_12 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__clkinv_12 I ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__aoi221_4 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__aoi221_4 A1 A2 B1 B2 C ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__nand3_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__nand3_2 A1 A2 A3 ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__and2_4 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__and2_4 A1 A2 Z VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__tieh abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__tieh Z VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 I Z VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__and4_4 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__and4_4 A1 A2 A3 A4 Z VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__mux2_4 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__mux2_4 I0 I1 S Z VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__inv_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__inv_1 I ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__and3_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__and3_2 A1 A2 A3 Z VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__oai221_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__oai221_2 A1 A2 B1 B2 C ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__aoi22_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__aoi22_2 A1 A2 B1 B2 ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__oai221_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__oai221_1 A1 A2 B1 B2 C ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__inv_3 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__inv_3 I ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__clkbuf_8 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__clkbuf_8 I Z VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__aoi21_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__aoi21_2 A1 A2 B ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__buf_3 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__buf_3 I Z VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__xnor2_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__xnor2_1 A1 A2 ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__oai22_4 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__oai22_4 A1 A2 B1 B2 ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__or4_4 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__or4_4 A1 A2 A3 A4 Z VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__aoi221_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__aoi221_2 A1 A2 B1 B2 C ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__buf_20 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__buf_20 I Z VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__buf_16 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__buf_16 I Z VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__and2_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__and2_2 A1 A2 Z VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__oai211_4 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__oai211_4 A1 A2 B C ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 I Z VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__and4_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__and4_2 A1 A2 A3 A4 Z VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__clkinv_8 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__clkinv_8 I ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__clkinv_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__clkinv_2 I ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__buf_8 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__buf_8 I Z VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__inv_8 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__inv_8 I ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__oai33_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__oai33_1 A1 A2 A3 B1 B2 B3 ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__inv_4 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__inv_4 I ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__aoi22_4 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__aoi22_4 A1 A2 B1 B2 ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__aoi222_4 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__aoi222_4 A1 A2 B1 B2 C1 C2 ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__oai22_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__oai22_2 A1 A2 B1 B2 ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__xor2_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__xor2_2 A1 A2 Z VDD VSS
.ends

.subckt housekeeping VDD VSS debug_in debug_mode debug_oeb debug_out irq[0] irq[1]
+ irq[2] mask_rev_in[0] mask_rev_in[10] mask_rev_in[11] mask_rev_in[12] mask_rev_in[13]
+ mask_rev_in[14] mask_rev_in[15] mask_rev_in[16] mask_rev_in[17] mask_rev_in[18]
+ mask_rev_in[19] mask_rev_in[1] mask_rev_in[20] mask_rev_in[21] mask_rev_in[22] mask_rev_in[23]
+ mask_rev_in[24] mask_rev_in[25] mask_rev_in[26] mask_rev_in[27] mask_rev_in[28]
+ mask_rev_in[29] mask_rev_in[2] mask_rev_in[30] mask_rev_in[31] mask_rev_in[3] mask_rev_in[4]
+ mask_rev_in[5] mask_rev_in[6] mask_rev_in[7] mask_rev_in[8] mask_rev_in[9] mgmt_gpio_in[0]
+ mgmt_gpio_in[10] mgmt_gpio_in[11] mgmt_gpio_in[12] mgmt_gpio_in[13] mgmt_gpio_in[14]
+ mgmt_gpio_in[15] mgmt_gpio_in[16] mgmt_gpio_in[17] mgmt_gpio_in[18] mgmt_gpio_in[19]
+ mgmt_gpio_in[1] mgmt_gpio_in[20] mgmt_gpio_in[21] mgmt_gpio_in[22] mgmt_gpio_in[23]
+ mgmt_gpio_in[24] mgmt_gpio_in[25] mgmt_gpio_in[26] mgmt_gpio_in[27] mgmt_gpio_in[28]
+ mgmt_gpio_in[29] mgmt_gpio_in[2] mgmt_gpio_in[30] mgmt_gpio_in[31] mgmt_gpio_in[32]
+ mgmt_gpio_in[33] mgmt_gpio_in[34] mgmt_gpio_in[35] mgmt_gpio_in[36] mgmt_gpio_in[37]
+ mgmt_gpio_in[3] mgmt_gpio_in[4] mgmt_gpio_in[5] mgmt_gpio_in[6] mgmt_gpio_in[7]
+ mgmt_gpio_in[8] mgmt_gpio_in[9] mgmt_gpio_oeb[0] mgmt_gpio_oeb[10] mgmt_gpio_oeb[11]
+ mgmt_gpio_oeb[12] mgmt_gpio_oeb[13] mgmt_gpio_oeb[14] mgmt_gpio_oeb[15] mgmt_gpio_oeb[16]
+ mgmt_gpio_oeb[17] mgmt_gpio_oeb[18] mgmt_gpio_oeb[19] mgmt_gpio_oeb[1] mgmt_gpio_oeb[20]
+ mgmt_gpio_oeb[21] mgmt_gpio_oeb[22] mgmt_gpio_oeb[23] mgmt_gpio_oeb[24] mgmt_gpio_oeb[25]
+ mgmt_gpio_oeb[26] mgmt_gpio_oeb[27] mgmt_gpio_oeb[28] mgmt_gpio_oeb[29] mgmt_gpio_oeb[2]
+ mgmt_gpio_oeb[30] mgmt_gpio_oeb[31] mgmt_gpio_oeb[32] mgmt_gpio_oeb[33] mgmt_gpio_oeb[34]
+ mgmt_gpio_oeb[35] mgmt_gpio_oeb[36] mgmt_gpio_oeb[37] mgmt_gpio_oeb[3] mgmt_gpio_oeb[4]
+ mgmt_gpio_oeb[5] mgmt_gpio_oeb[6] mgmt_gpio_oeb[7] mgmt_gpio_oeb[8] mgmt_gpio_oeb[9]
+ mgmt_gpio_out[0] mgmt_gpio_out[10] mgmt_gpio_out[11] mgmt_gpio_out[12] mgmt_gpio_out[13]
+ mgmt_gpio_out[14] mgmt_gpio_out[15] mgmt_gpio_out[16] mgmt_gpio_out[17] mgmt_gpio_out[18]
+ mgmt_gpio_out[19] mgmt_gpio_out[1] mgmt_gpio_out[20] mgmt_gpio_out[21] mgmt_gpio_out[22]
+ mgmt_gpio_out[23] mgmt_gpio_out[24] mgmt_gpio_out[25] mgmt_gpio_out[26] mgmt_gpio_out[27]
+ mgmt_gpio_out[28] mgmt_gpio_out[29] mgmt_gpio_out[2] mgmt_gpio_out[30] mgmt_gpio_out[31]
+ mgmt_gpio_out[32] mgmt_gpio_out[33] mgmt_gpio_out[34] mgmt_gpio_out[35] mgmt_gpio_out[36]
+ mgmt_gpio_out[37] mgmt_gpio_out[3] mgmt_gpio_out[4] mgmt_gpio_out[5] mgmt_gpio_out[6]
+ mgmt_gpio_out[7] mgmt_gpio_out[8] mgmt_gpio_out[9] pad_flash_clk pad_flash_clk_oe
+ pad_flash_csb pad_flash_csb_oe pad_flash_io0_di pad_flash_io0_do pad_flash_io0_ie
+ pad_flash_io0_oe pad_flash_io1_di pad_flash_io1_do pad_flash_io1_ie pad_flash_io1_oe
+ pll90_sel[0] pll90_sel[1] pll90_sel[2] pll_bypass pll_dco_ena pll_div[0] pll_div[1]
+ pll_div[2] pll_div[3] pll_div[4] pll_ena pll_sel[0] pll_sel[1] pll_sel[2] pll_trim[0]
+ pll_trim[10] pll_trim[11] pll_trim[12] pll_trim[13] pll_trim[14] pll_trim[15] pll_trim[16]
+ pll_trim[17] pll_trim[18] pll_trim[19] pll_trim[1] pll_trim[20] pll_trim[21] pll_trim[22]
+ pll_trim[23] pll_trim[24] pll_trim[25] pll_trim[2] pll_trim[3] pll_trim[4] pll_trim[5]
+ pll_trim[6] pll_trim[7] pll_trim[8] pll_trim[9] porb pwr_ctrl_out qspi_enabled reset
+ ser_rx ser_tx serial_clock serial_data_1 serial_data_2 serial_load serial_resetn
+ spi_csb spi_enabled spi_sck spi_sdi spi_sdo spi_sdoenb spimemio_flash_clk spimemio_flash_csb
+ spimemio_flash_io0_di spimemio_flash_io0_do spimemio_flash_io0_oeb spimemio_flash_io1_di
+ spimemio_flash_io1_do spimemio_flash_io1_oeb spimemio_flash_io2_di spimemio_flash_io2_do
+ spimemio_flash_io2_oeb spimemio_flash_io3_di spimemio_flash_io3_do spimemio_flash_io3_oeb
+ trap uart_enabled user_clock wb_ack_o wb_adr_i[0] wb_adr_i[10] wb_adr_i[11] wb_adr_i[12]
+ wb_adr_i[13] wb_adr_i[14] wb_adr_i[15] wb_adr_i[16] wb_adr_i[17] wb_adr_i[18] wb_adr_i[19]
+ wb_adr_i[1] wb_adr_i[20] wb_adr_i[21] wb_adr_i[22] wb_adr_i[23] wb_adr_i[24] wb_adr_i[25]
+ wb_adr_i[26] wb_adr_i[27] wb_adr_i[28] wb_adr_i[29] wb_adr_i[2] wb_adr_i[30] wb_adr_i[31]
+ wb_adr_i[3] wb_adr_i[4] wb_adr_i[5] wb_adr_i[6] wb_adr_i[7] wb_adr_i[8] wb_adr_i[9]
+ wb_clk_i wb_cyc_i wb_dat_i[0] wb_dat_i[10] wb_dat_i[11] wb_dat_i[12] wb_dat_i[13]
+ wb_dat_i[14] wb_dat_i[15] wb_dat_i[16] wb_dat_i[17] wb_dat_i[18] wb_dat_i[19] wb_dat_i[1]
+ wb_dat_i[20] wb_dat_i[21] wb_dat_i[22] wb_dat_i[23] wb_dat_i[24] wb_dat_i[25] wb_dat_i[26]
+ wb_dat_i[27] wb_dat_i[28] wb_dat_i[29] wb_dat_i[2] wb_dat_i[30] wb_dat_i[31] wb_dat_i[3]
+ wb_dat_i[4] wb_dat_i[5] wb_dat_i[6] wb_dat_i[7] wb_dat_i[8] wb_dat_i[9] wb_dat_o[0]
+ wb_dat_o[10] wb_dat_o[11] wb_dat_o[12] wb_dat_o[13] wb_dat_o[14] wb_dat_o[15] wb_dat_o[16]
+ wb_dat_o[17] wb_dat_o[18] wb_dat_o[19] wb_dat_o[1] wb_dat_o[20] wb_dat_o[21] wb_dat_o[22]
+ wb_dat_o[23] wb_dat_o[24] wb_dat_o[25] wb_dat_o[26] wb_dat_o[27] wb_dat_o[28] wb_dat_o[29]
+ wb_dat_o[2] wb_dat_o[30] wb_dat_o[31] wb_dat_o[3] wb_dat_o[4] wb_dat_o[5] wb_dat_o[6]
+ wb_dat_o[7] wb_dat_o[8] wb_dat_o[9] wb_rstn_i wb_sel_i[0] wb_sel_i[1] wb_sel_i[2]
+ wb_sel_i[3] wb_stb_i wb_we_i
XFILLER_100_138 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_67_553 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_39_211 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_54_203 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_55_726 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_7963_ _7963_/D _7316_/Z _7972_/CLK _7963_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffnsnq_1
XFILLER_94_372 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_82_534 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_67_597 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_27_428 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_82_567 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6914_ _6955_/A4 _6935_/A2 _7202_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_4
XFILLER_54_247 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_54_258 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_35_461 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7894_ _7894_/D _7900_/RN _7900_/CLK _7894_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffsnq_1
X_6845_ _7667_/Q _6885_/A2 _6647_/Z _7619_/Q _6887_/B1 _7683_/Q _6847_/A2 VDD VSS
+ gf180mcu_fd_sc_mcu7t5v0__aoi222_1
XFILLER_168_18 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3988_ _7625_/Q _5954_/A1 _6226_/A1 _7753_/Q _3989_/A4 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_6776_ _6776_/A1 _6776_/A2 _6776_/A3 _6776_/A4 _6777_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand4_1
X_5727_ _5331_/Z _5727_/A2 _5437_/B _5619_/Z _5763_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand4_2
XFILLER_176_694 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_164_812 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_175_171 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_148_396 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5658_ _5669_/A1 _5179_/B _5658_/B _5674_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_5589_ _5589_/A1 _5589_/A2 _5589_/A3 _5590_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor3_1
X_4609_ _4609_/A1 _6537_/A2 _4613_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_7328_ _7901_/RN _4334_/Z _7328_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_144_591 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_117_783 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_116_271 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xhold340 _7609_/Q hold340/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
Xhold351 hold351/I _6204_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
Xhold362 hold362/I _7362_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
X_7259_ _7518_/Q _7259_/A2 _7261_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
Xhold373 hold373/I _6328_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
XFILLER_89_144 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
Xhold384 _7624_/Q hold384/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
Xhold395 hold395/I _7537_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
XFILLER_131_274 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_117_99 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_131_296 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_58_520 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_58_542 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_100_672 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_85_372 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1800 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_93_58 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_73_567 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_165_2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1833 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1822 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1811 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_159_617 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1866 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1855 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1844 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_158_127 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_158_105 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1899 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1888 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1877 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_13_144 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_167_650 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_155_812 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_166_193 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_127_558 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_182_664 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_181_141 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_170_804 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_5_354 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_123_753 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_68_328 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_110_458 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_110_447 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_49_531 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_67_70 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_64_534 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_36_203 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_36_247 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4960_ _5797_/B _4965_/B _4960_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__or2_1
XFILLER_45_770 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_3911_ _3911_/A1 _3911_/A2 _3911_/A3 _3911_/A4 _3917_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand4_1
X_4891_ hold850/Z _4892_/A2 _4892_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_177_425 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_149_127 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3842_ hold72/I hold54/Z hold55/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_4
X_6630_ _7907_/Q _6633_/A2 _6664_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_4
XFILLER_80_2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6561_ _7902_/Q _7903_/Q _6561_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_164_108 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3773_ _4292_/B _3774_/A2 _7965_/Q _3774_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_146_812 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5512_ _5621_/B _5648_/B2 _5512_/B _5514_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_173_631 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6492_ _4460_/Z _6502_/A2 _6492_/B _7872_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_9_682 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5443_ _5621_/B _5648_/B2 _5629_/B _5572_/B _5444_/A4 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XFILLER_160_325 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5374_ _5405_/B _5504_/A3 _5577_/B2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_4325_ _4309_/S _4325_/A2 _4325_/B _7336_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_113_241 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_7113_ _7796_/Q _7190_/A2 _7190_/B1 _7618_/Q _7190_/C1 _7706_/Q _7116_/A2 VDD VSS
+ gf180mcu_fd_sc_mcu7t5v0__aoi222_1
XFILLER_101_425 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7044_ _7623_/Q _7195_/B1 _7200_/B1 hold98/I _7048_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_4256_ _4256_/A1 _4256_/A2 _4256_/A3 _4256_/A4 _4263_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand4_1
X_4187_ _4187_/A1 _4187_/A2 _4187_/A3 _4187_/A4 _4203_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor4_2
XFILLER_95_692 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_55_523 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_55_567 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1118 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1129 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_7946_ _7946_/D _7949_/CLK _7946_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_1107 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_228 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_7877_ _7877_/D _7877_/RN _7877_/CLK _7877_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_70_559 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_6828_ _7927_/Q _7133_/S _6829_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_50_250 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_137_6 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_11_637 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_137_812 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6759_ _7728_/Q _6892_/B1 _6880_/B1 _7810_/Q _6766_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_163_141 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_128_54 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_151_303 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_128_65 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_117_580 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_105_753 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xhold170 _7889_/Q hold170/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
Xhold192 _7339_/Q hold192/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
XFILLER_78_637 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_2_379 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xhold181 hold181/I _7639_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
XFILLER_144_64 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_120_756 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_144_86 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_46_534 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_58_383 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2320 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_18_247 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_37_73 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_2353 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2342 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2331 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2386 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2375 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2364 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1641 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1630 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2397 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_159_425 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1685 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1674 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1663 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1652 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1696 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_146_119 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_146_108 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_128_812 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_127_377 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_142_347 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_142_336 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_111_701 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_111_712 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_123_583 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5090_ _5692_/B _5285_/A3 _5424_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_2
X_4110_ _4110_/I0 hold947/Z _4427_/B _7550_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_4041_ _7719_/Q hold90/I _4046_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_96_467 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_68_158 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_68_169 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_49_372 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_37_567 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_92_673 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7800_ _7800_/D _7901_/RN _7901_/CLK _7800_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffsnq_1
X_5992_ _4454_/Z _6004_/A2 _5992_/B _7637_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_37_578 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4943_ _3728_/I _4900_/Z _4943_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__xor2_4
X_7731_ _7731_/D _7877_/RN _7852_/CLK _7731_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_33_740 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_7662_ _7662_/D _7877_/RN _7849_/CLK _7662_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffsnq_1
XFILLER_32_250 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6613_ _7915_/Q _6905_/A2 _6955_/A4 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_4
X_4874_ hold604/Z _4877_/A2 hold605/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_165_428 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_119_812 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3825_ hold38/Z _4212_/A2 _6056_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_4
X_7593_ _7593_/D _7900_/RN _7892_/CLK _8003_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
X_3756_ _4383_/A2 _3772_/S _4291_/A2 _3756_/B _3765_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai31_2
X_6544_ hold176/Z _6553_/A2 hold177/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_20_478 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_145_141 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6475_ _4460_/Z _6485_/A2 _6475_/B _7864_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_3687_ _7801_/Q _3687_/ZN VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_5426_ _5712_/B _5534_/A2 _5691_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_161_645 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
Xoutput242 _7986_/Z mgmt_gpio_out[5] VDD VSS gf180mcu_fd_sc_mcu7t5v0__buf_4
Xoutput253 _4422_/I pad_flash_io0_oe VDD VSS gf180mcu_fd_sc_mcu7t5v0__buf_4
Xoutput220 _4404_/ZN mgmt_gpio_out[1] VDD VSS gf180mcu_fd_sc_mcu7t5v0__buf_4
Xoutput231 _7983_/Z mgmt_gpio_out[2] VDD VSS gf180mcu_fd_sc_mcu7t5v0__buf_4
X_5357_ _5357_/A1 _5643_/A2 _5667_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_114_550 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xoutput286 _7354_/Q pll_trim[23] VDD VSS gf180mcu_fd_sc_mcu7t5v0__buf_4
Xoutput264 _7560_/Q pll_div[2] VDD VSS gf180mcu_fd_sc_mcu7t5v0__buf_4
Xoutput275 _7360_/Q pll_trim[13] VDD VSS gf180mcu_fd_sc_mcu7t5v0__buf_4
XFILLER_181_18 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4308_ _3808_/Z _4308_/I1 _4308_/S _4308_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_99_283 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5288_ _5288_/A1 _5288_/A2 _5288_/A3 _5288_/A4 _5298_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand4_1
XFILLER_87_445 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xoutput297 _7572_/Q pwr_ctrl_out VDD VSS gf180mcu_fd_sc_mcu7t5v0__buf_4
XFILLER_114_23 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_101_266 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7027_ _7027_/A1 _7210_/A2 _7027_/B _7433_/Q _7028_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi211_1
X_4239_ input20/Z _4239_/A2 _4774_/A1 _7474_/Q _4240_/A4 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_28_534 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7929_ _7929_/D _7938_/RN _7940_/CLK _7929_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_169_712 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_90_37 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_11_423 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_23_261 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_24_784 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_51_570 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_128_108 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_11_434 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_128_2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_7_416 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_99_68 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_99_57 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_3_611 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_151_144 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_2_121 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_151_166 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_112_509 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_120_531 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_120_520 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_2_176 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_120_575 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_78_489 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_171_73 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_68 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_46 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_19_567 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2161 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2150 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2194 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2183 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2172 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1460 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1493 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1482 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1471 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_14_250 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_9_33 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_147_428 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_80_70 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4590_ hold754/Z _4593_/A2 _4591_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_127_141 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_127_130 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_155_483 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_143_623 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
Xhold906 hold906/I _7557_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
XFILLER_6_460 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xhold928 _7741_/Q hold928/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
Xhold917 hold917/I _6196_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
Xhold939 _7955_/Q _3672_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
X_6260_ _6549_/A1 _6264_/A2 _6260_/B _7763_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_5211_ _3723_/I _4906_/S _5211_/A3 _4920_/Z _5373_/A4 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand4_4
X_6191_ _6553_/A1 _6191_/A2 _6191_/B _7731_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_103_509 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_43_2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5142_ _5309_/A1 _3723_/I _5006_/B _5254_/A2 _5545_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand4_4
XFILLER_29_309 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5073_ _4943_/Z _4993_/B _5663_/A1 _5077_/C VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor3_1
X_4024_ _4024_/A1 _4024_/A2 _4024_/A3 _4024_/A4 _4025_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand4_1
XFILLER_49_191 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_92_481 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_25_548 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5975_ _4454_/Z _5987_/A2 _5975_/B _7629_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_80_676 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_178_531 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4926_ _4926_/A1 _4926_/A2 _4926_/A3 _4926_/A4 _4926_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__or4_2
X_7714_ _7714_/D _7853_/RN _7811_/CLK _7714_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_33_570 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_52_389 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_178_575 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4857_ _4454_/Z _4857_/A2 _4857_/B hold811/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_7645_ _7645_/D _7961_/RN _7649_/CLK _7645_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffsnq_1
X_3808_ hold147/Z hold192/Z _7414_/Q _3808_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_7576_ hold65/Z _7961_/RN _7624_/CLK _7576_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_181_729 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_6527_ hold170/Z _6536_/A2 hold171/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_4788_ _7221_/A1 _4795_/S _4788_/B _7479_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_174_770 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3739_ _7344_/Q _3730_/Z _4383_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_118_185 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_106_325 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6458_ _4460_/Z _6468_/A2 _6458_/B _7856_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_133_177 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_133_144 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5409_ _4993_/C _5099_/B _5645_/A3 _5409_/B2 _5411_/C VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai22_1
X_6389_ hold686/Z _6400_/A2 _6390_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_121_339 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_102_531 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_614 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_125_55 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_87_286 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_28_342 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_56_684 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_83_481 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_70_120 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_70_175 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_24_581 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_34_41 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_12_732 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_24_592 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_129_428 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_8_747 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_156_269 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_156_247 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_11_286 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_7_224 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_7_235 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_50_62 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_164_280 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_152_442 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_152_475 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_125_667 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_507 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_78_220 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_529 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_518 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_3_496 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_3_485 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_182_72 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_120_372 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_93_212 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_93_267 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_75_70 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_34_301 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_62_676 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5760_ _5617_/Z _5684_/Z _5760_/A3 _5760_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__and3_1
XFILLER_15_570 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_22_529 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_34_389 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4711_ _7442_/Q _4718_/A1 _4714_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_5691_ _5691_/A1 _5622_/Z _5691_/A3 _5691_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__and3_1
XTAP_1290 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_7430_ _7430_/D _7853_/RN _7601_/CLK _7430_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
X_4642_ _3830_/Z _4476_/I _4643_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_175_567 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xhold703 hold703/I _7698_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
X_7361_ _7361_/D _7875_/RN _7410_/CLK _7361_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffsnq_1
X_4573_ _4454_/Z _4573_/A2 _4573_/B _7392_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_7292_ _7901_/RN _4334_/Z _7292_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__and2_1
Xhold725 _7787_/Q hold725/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
X_6312_ hold307/Z _6315_/A2 _6313_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
Xhold714 hold714/I _7682_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
XFILLER_7_780 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xhold736 hold736/I _4880_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
XFILLER_170_250 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_143_453 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_115_144 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xhold747 hold747/I _7360_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
Xhold769 _7397_/Q hold769/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
X_6243_ _6243_/A1 _6537_/A2 _6247_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
Xhold758 _7677_/Q hold758/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
XFILLER_131_659 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_131_626 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_130_125 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_130_103 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6174_ _6553_/A1 _6174_/A2 _6174_/B hold156/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_5125_ _5543_/C _5543_/B _5479_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_69_286 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_29_106 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5056_ _5199_/B _3727_/I _3728_/I _5369_/B _5087_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor4_4
XFILLER_85_779 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_84_234 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_84_256 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4007_ hold76/Z hold149/Z _5817_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_4
XFILLER_65_492 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_38_695 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_80_495 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5958_ _4454_/Z _5970_/A2 _5958_/B _7621_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_4909_ _4925_/A1 _4923_/A1 _4914_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_21_540 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_52_197 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_166_534 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_5889_ hold826/Z _5902_/A2 _5890_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_7628_ _7628_/D _7877_/RN _7809_/CLK _7628_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffsnq_1
XFILLER_138_247 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_153_228 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_7559_ _7559_/D _7875_/RN _7563_/CLK _7559_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_147_792 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_161_283 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_422 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xhold30 hold30/I hold30/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
Xhold41 hold41/I hold41/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
XFILLER_76_735 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_75_212 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_48_404 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xhold63 hold63/I hold63/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
XFILLER_152_64 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
Xhold74 hold74/I hold74/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
Xhold52 hold52/I hold52/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
XFILLER_75_223 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_48_437 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_152_86 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
Xhold85 hold85/I hold85/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
Xhold96 hold96/I hold96/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
XFILLER_28_183 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_44_632 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xclkbuf_3_7__f_wb_clk_i clkbuf_0_wb_clk_i/Z _4411_/I1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_28_194 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_43_131 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_45_73 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_44_676 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_351 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_340 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_362 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_169_383 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_129_225 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_8_500 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_157_567 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_172_504 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_157_578 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_8_577 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_152_250 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_152_283 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_152_261 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_140_401 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_112_103 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_3_293 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_100_309 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_39_404 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_39_459 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_67_779 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_66_256 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_54_407 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_54_418 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_81_215 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6930_ _7914_/Q _7913_/Q _6599_/Z _6941_/A2 _7190_/B1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor4_4
Xclkbuf_leaf_6_csclk clkbuf_leaf_9_csclk/I _7898_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
X_6861_ _7399_/Q _6894_/A2 _6891_/A2 _7407_/Q _6864_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_6792_ _7689_/Q _6884_/B1 _6792_/B _6792_/C _6800_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XFILLER_62_473 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_5812_ _5812_/A1 _6537_/A2 _5816_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_50_602 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5743_ _5743_/A1 _5743_/A2 _5743_/A3 _5766_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_50_635 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_176_810 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_148_534 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5674_ _5674_/A1 _5674_/A2 _5674_/A3 _5773_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_30_392 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4625_ _7991_/I _4652_/A1 _4628_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_7413_ _7413_/D _7304_/Z _4415_/A2 _7413_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_2
XFILLER_163_526 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_129_770 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7344_ _7344_/D _7299_/Z _4398_/I1 _7344_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_2
XFILLER_128_291 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
Xhold511 hold511/I _6070_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
Xhold500 _7604_/Q hold500/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
X_4556_ _6539_/A1 _4558_/A2 _4556_/B _7385_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
Xhold522 hold522/I _7430_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
Xhold544 hold544/I _7680_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
Xhold533 _7874_/Q hold533/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
Xhold566 hold566/I _7416_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
X_7275_ _7520_/Q _7275_/A2 _7275_/B1 _7519_/Q _7276_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_171_570 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xhold577 hold577/I _7710_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
XFILLER_143_283 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_131_401 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_116_475 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
Xhold588 _7762_/Q hold588/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
Xhold555 hold555/I _6202_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
X_4487_ _4487_/A1 _6553_/A1 _4487_/B _7354_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_6226_ _6226_/A1 _7285_/A2 hold6/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_4
Xhold599 hold599/I _7523_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
X_6157_ _6553_/A1 _6157_/A2 _6157_/B hold304/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_131_489 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_106_57 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_860 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_871 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_58_724 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5108_ _5661_/A1 _5797_/C _5647_/A2 _5672_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor3_4
XFILLER_97_392 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_882 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_893 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_57_212 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6088_ hold184/Z _6089_/A2 hold185/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_5039_ _5151_/A1 _5151_/A2 _5041_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_122_34 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_26_654 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_13_304 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_25_175 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_26_676 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_41_602 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_167_810 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_139_545 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_5_514 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_110_2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_134_250 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_181_389 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_134_283 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_1_753 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
Xinput120 wb_adr_i[3] _5006_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__buf_12
XFILLER_0_263 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
Xinput142 wb_dat_i[22] _7270_/B1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyb_1
Xinput153 wb_dat_i[3] _7257_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyb_1
Xinput131 wb_dat_i[12] _7260_/B1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XFILLER_88_392 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xinput164 wb_sel_i[3] _7281_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XFILLER_63_226 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_63_215 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_44_440 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_44_495 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_177_629 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_170 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_32_668 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_192 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_181 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_31_189 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_157_386 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_12_392 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_172_312 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4410_ _7443_/Q user_clock _7584_/Q _4410_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_68_4 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_160_518 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5390_ _5660_/A2 _5390_/A2 _5701_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_99_602 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_172_389 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4341_ _7519_/Q _4438_/A2 _7514_/Q _4342_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_160_529 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_153_570 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_125_283 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_98_101 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_98_156 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_7060_ _7802_/Q _7191_/B1 _7190_/C1 _7704_/Q _7063_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_4272_ _7363_/Q _4505_/A1 _4569_/A1 _7391_/Q _4274_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_6011_ _4460_/Z _6021_/A2 _6011_/B _7646_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_79_392 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7962_ _7962_/D _7315_/Z _4415_/A2 hold21/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffnrnq_1
X_6913_ _7914_/Q _7913_/Q _6936_/A1 _6935_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand3_4
X_7893_ _7893_/D _7901_/RN _7899_/CLK _7893_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
X_6844_ _7805_/Q _6883_/A2 _6883_/B1 _7789_/Q _6884_/B1 _7691_/Q _6847_/A1 VDD VSS
+ gf180mcu_fd_sc_mcu7t5v0__aoi222_1
XFILLER_167_106 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3987_ _7705_/Q _6124_/A1 _6107_/A1 _7697_/Q _3989_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_6775_ _7712_/Q _6885_/B1 _6890_/A2 _7640_/Q _6776_/A4 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_5726_ _5726_/A1 _5726_/A2 _5761_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_10_318 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_182_109 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_176_673 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_175_150 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_109_707 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5657_ _5706_/A1 _5657_/A2 _5657_/A3 _5657_/A4 _5657_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__and4_1
X_5588_ _5673_/A2 _5566_/B _5588_/A3 _5733_/A3 _5589_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand4_1
X_4608_ _4454_/Z _4608_/A2 _4608_/B _7406_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_4539_ hold183/Z _4548_/A2 _4540_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_7327_ _7901_/RN _4334_/Z _7327_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__and2_1
Xhold330 hold330/I _6119_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
XFILLER_117_45 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_116_250 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
Xhold341 hold341/I _5932_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
Xhold352 hold352/I _7737_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
X_7258_ _7258_/A1 _7277_/B _7258_/B _7953_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi21_1
Xhold374 hold374/I _7795_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
XFILLER_117_56 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
Xhold363 _7676_/Q hold363/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
Xhold385 _7575_/Q hold385/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
Xhold396 _7648_/Q hold396/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
XFILLER_104_478 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_104_489 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_6209_ hold43/Z hold5/Z _6225_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_4
XFILLER_131_286 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_7189_ _7528_/Q _7189_/A2 _7189_/B1 _7522_/Q _7189_/C1 _7495_/Q _7192_/A1 VDD VSS
+ gf180mcu_fd_sc_mcu7t5v0__aoi222_1
XTAP_690 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_18_429 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_45_215 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_61_708 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1834 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1823 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1812 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1801 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_54_760 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_158_2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1867 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1856 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1845 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_14_646 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_41_432 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_53_281 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1889 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1878 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_158_52 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_6_812 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_182_632 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_154_334 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_5_344 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_154_389 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_135_570 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_123_765 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_107_283 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_69_808 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_122_275 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_96_616 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_96_605 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_68_318 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_92_811 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_67_82 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
Xclkbuf_leaf_71_csclk clkbuf_3_3__f_csclk/Z _7639_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_91_354 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_83_70 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3910_ _7739_/Q _6192_/A1 _6107_/A1 _7699_/Q _3911_/A4 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_1
Xclkbuf_leaf_86_csclk _7528_/CLK _7401_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
X_4890_ _6539_/A1 _4892_/A2 _4890_/B _7535_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_149_106 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3841_ _4212_/A2 _4141_/A1 _6192_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_4
XFILLER_20_605 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3772_ input58/Z hold967/Z _3772_/S _7966_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_32_498 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6560_ _7902_/Q _6564_/B _6560_/B _7902_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_158_673 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5511_ _5648_/A1 _5669_/B _5431_/B _5648_/B2 _5511_/C _5514_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi221_1
XFILLER_118_515 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_118_504 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_73_2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_158_695 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_157_172 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6491_ hold696/Z _6502_/A2 _6492_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_5442_ _5319_/C _5563_/B2 _5687_/B _5319_/B _5692_/A2 _5629_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai32_1
XFILLER_8_193 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_173_698 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_5373_ _4906_/Z _5585_/A1 _5373_/A3 _5373_/A4 _5576_/B2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand4_2
X_4324_ _7336_/Q _4309_/S _4325_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
Xclkbuf_leaf_24_csclk _7422_/CLK _7849_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
X_7112_ _7682_/Q _7191_/A2 _7116_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_7043_ _7043_/A1 _7043_/A2 _7043_/A3 _7054_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_113_286 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_87_638 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4255_ _7748_/Q _6226_/A1 _6243_/A1 _7756_/Q _4256_/A4 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_1
Xclkbuf_leaf_39_csclk clkbuf_3_7__f_csclk/Z _7755_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_83_800 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_67_351 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4186_ _4186_/A1 _4186_/A2 _4187_/A4 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_95_682 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_27_215 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_55_535 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_82_321 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_27_237 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_55_546 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_7945_ _7945_/D _7949_/CLK _7945_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_1119 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1108 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_23_432 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_35_292 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7876_ _7876_/D _7961_/RN _7876_/CLK _7876_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
X_6827_ _7433_/Q _7926_/Q _6827_/B _6829_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_168_437 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6758_ _7794_/Q _6893_/A2 _6890_/B1 hold59/I _6766_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_6_108 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_164_632 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5709_ _5709_/A1 _5709_/A2 _5710_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_6689_ _7791_/Q _6893_/A2 _6893_/B1 _7767_/Q _6692_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_164_676 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_124_507 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_136_389 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_124_529 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_117_570 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_88_37 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_128_99 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_117_592 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xhold160 _7857_/Q hold160/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
Xhold171 hold171/I _6528_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
Xhold193 _3781_/Z hold193/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
Xhold182 _7833_/Q hold182/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
XFILLER_78_605 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_19_705 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_74_811 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_19_749 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_2310 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2343 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2332 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2321 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_73_354 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2387 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2376 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2354 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2365 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_160_97 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1642 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1631 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1620 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2398 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_159_415 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1675 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1664 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1653 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_763 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1697 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1686 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_53_73 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_169_73 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_127_312 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_182_440 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_170_602 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_10_682 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_6_664 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_5_141 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_170_646 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_150_392 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_110_212 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_69_638 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4040_ _7889_/Q _6520_/A1 _4719_/A1 input64/Z _4052_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_65_800 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_64_321 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5991_ hold884/Z _6004_/A2 _5992_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_4942_ _4920_/Z _4973_/A3 _4942_/B _5600_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_4
X_7730_ _7730_/D _7877_/RN _7852_/CLK _7730_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_64_387 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_178_735 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_177_212 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7661_ _7661_/D _7877_/RN _7849_/CLK _7661_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffsnq_1
X_6612_ _6612_/I _7915_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_4873_ _4873_/A1 _7285_/A2 _4877_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_3824_ _3783_/Z hold41/Z hold75/Z _3963_/A4 _4212_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand4_4
XFILLER_20_435 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7592_ _7592_/D _7900_/RN _7592_/CLK _8002_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
X_3755_ _7413_/Q _3738_/Z _4291_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_6543_ _4460_/Z _6553_/A2 _6543_/B hold592/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_3686_ _7809_/Q _3686_/ZN VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_6474_ hold669/Z _6485_/A2 _6475_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_161_635 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_146_676 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_145_153 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_118_389 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5425_ _5062_/Z _5176_/B _5425_/B _5437_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_2
Xoutput210 _4397_/Z mgmt_gpio_out[10] VDD VSS gf180mcu_fd_sc_mcu7t5v0__buf_4
XFILLER_160_112 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
Xoutput232 _8004_/Z mgmt_gpio_out[30] VDD VSS gf180mcu_fd_sc_mcu7t5v0__buf_4
XFILLER_133_359 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xoutput221 _7994_/Z mgmt_gpio_out[20] VDD VSS gf180mcu_fd_sc_mcu7t5v0__buf_4
Xoutput243 _4400_/Z mgmt_gpio_out[6] VDD VSS gf180mcu_fd_sc_mcu7t5v0__buf_4
X_5356_ _5094_/C _5356_/A2 _5356_/A3 _5356_/A4 _5359_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand4_1
Xoutput254 _8007_/Z pad_flash_io1_do VDD VSS gf180mcu_fd_sc_mcu7t5v0__buf_4
Xoutput276 _7361_/Q pll_trim[14] VDD VSS gf180mcu_fd_sc_mcu7t5v0__buf_4
XFILLER_0_807 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xoutput265 _7561_/Q pll_div[3] VDD VSS gf180mcu_fd_sc_mcu7t5v0__buf_4
X_4307_ _4306_/Z _7341_/Q _4309_/S _7341_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_141_370 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5287_ _5575_/A2 _5425_/B _5287_/B _5287_/C _5288_/A4 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XFILLER_101_212 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xoutput298 _4215_/Z reset VDD VSS gf180mcu_fd_sc_mcu7t5v0__buf_4
Xoutput287 _7569_/Q pll_trim[24] VDD VSS gf180mcu_fd_sc_mcu7t5v0__buf_4
X_7026_ _7210_/A2 _7026_/A2 _7026_/A3 _7026_/A4 _7027_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor4_1
X_4238_ _7920_/Q _5870_/A1 _4238_/B1 input93/Z _4240_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_114_79 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_83_641 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_74_17 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4169_ _7847_/Q _6435_/A1 _4249_/A2 input15/Z _5881_/A1 _7587_/Q _4170_/A3 VDD VSS
+ gf180mcu_fd_sc_mcu7t5v0__aoi222_1
XFILLER_55_343 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_55_354 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_130_34 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_24_730 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_7928_ _7928_/D _7938_/RN _7938_/CLK _7928_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_169_724 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_130_56 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_168_212 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7859_ _7859_/D _7901_/RN _7864_/CLK _7859_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_169_779 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_137_621 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_7_428 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_136_120 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_99_47 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_152_602 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_140_808 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_124_337 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_3_2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_120_510 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_132_392 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_48_95 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_74_652 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_46_321 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_74_685 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_73_162 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_2162 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2151 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2140 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_64_50 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2195 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2184 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2173 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1450 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_61_357 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_61_346 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_159_212 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1483 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1472 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1461 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_14_273 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1494 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_30_744 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_9_89 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_30_788 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_127_120 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_128_676 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_115_304 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
Xhold907 _7364_/Q hold907/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
XFILLER_6_472 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
Xhold918 hold918/I _7733_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
X_5210_ _5087_/C _4914_/Z _5210_/A3 _5210_/B _5373_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai31_2
Xhold929 _7528_/Q hold929/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
X_6190_ hold315/Z _6191_/A2 _6191_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_130_318 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5141_ _3722_/I _5087_/C _5394_/A1 _5006_/C _5176_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor4_4
XFILLER_36_2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5072_ _5476_/B _5689_/A1 _5072_/B _5072_/C _5106_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_111_565 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_96_276 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4023_ _7810_/Q _6350_/A1 _6226_/A1 hold57/I _4024_/A4 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_38_800 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_65_641 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_92_460 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_65_663 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_37_354 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_25_538 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5974_ hold894/Z _5987_/A2 _5975_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_7713_ _7713_/D _7877_/RN _7726_/CLK _7713_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
X_4925_ _4925_/A1 input96/Z _4926_/A4 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_100_37 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_4856_ hold809/Z _4857_/A2 hold810/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_7644_ _7644_/D _7961_/RN _7649_/CLK _7644_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffsnq_1
XFILLER_165_215 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3807_ _7340_/Q _4383_/A1 _4308_/I1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_21_799 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_7575_ _7575_/D _7961_/RN _7624_/CLK _7575_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_165_248 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_118_120 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6526_ _4460_/Z _6536_/A2 _6526_/B hold595/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_4787_ _7479_/Q _4795_/S _4788_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_3738_ _7344_/Q _3730_/Z _3738_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_146_473 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_134_602 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_109_35 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3669_ _7952_/Q _7253_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_161_432 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_134_646 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_109_68 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6457_ hold586/Z _6468_/A2 _6458_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_5408_ _5585_/A1 _5608_/B _5621_/B _5759_/A1 _5408_/C _5413_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi221_1
X_6388_ _4454_/Z _6400_/A2 _6388_/B _7823_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_5339_ _5200_/B _3727_/I _4915_/Z _5422_/B _5618_/B1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand4_4
XFILLER_88_744 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_114_392 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_659 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_125_89 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_88_788 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_85_38 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_75_405 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7009_ _7848_/Q _7193_/A2 _7193_/C1 _7726_/Q _7193_/B1 _7630_/Q _7016_/A1 VDD VSS
+ gf180mcu_fd_sc_mcu7t5v0__aoi222_1
XFILLER_87_298 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_28_332 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_28_321 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_141_44 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
Xclkbuf_3_6__f_wb_clk_i clkbuf_0_wb_clk_i/Z _7935_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_31_508 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_43_357 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_140_2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_12_744 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_11_210 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_156_259 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_137_495 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_109_186 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_140_605 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_79_700 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_112_318 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_112_329 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_519 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_508 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_105_392 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_79_777 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_78_254 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_94_747 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_47_641 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_75_82 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_19_354 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_61_132 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_34_335 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_61_154 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_34_379 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4710_ _4718_/A1 _4710_/A2 _4710_/B hold508/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_5690_ _5690_/A1 _5757_/A2 _5691_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_91_70 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1291 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1280 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_148_727 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_147_215 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4641_ hold692/Z _4652_/A1 _4644_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_147_248 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_30_585 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_30_596 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_116_602 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7360_ _7360_/D _7961_/RN _7570_/CLK _7360_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffsnq_1
X_4572_ hold851/Z _4573_/A2 _4573_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_7291_ _7901_/RN _4334_/Z _7291_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_155_292 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xhold726 _7763_/Q hold726/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
X_6311_ _6549_/A1 _6315_/A2 _6311_/B _7787_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
Xhold715 _7820_/Q hold715/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
Xhold737 hold737/I _7531_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
Xhold704 _7568_/Q hold704/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
X_6242_ hold2/Z hold6/Z _6242_/B hold7/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_115_167 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_104_808 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xhold748 _7756_/Q hold748/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
Xhold759 hold759/I _6077_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
XFILLER_131_638 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6173_ hold155/Z _6174_/A2 _6174_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_5124_ _5533_/A1 _5543_/B _5540_/B1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_5055_ _3728_/I _5369_/B _5421_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_4
X_4006_ _7858_/Q _6452_/A1 _4035_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_93_780 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_25_357 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_41_806 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_111_69 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_80_463 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_13_508 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5957_ hold881/Z _5970_/A2 _5958_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_52_176 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4908_ _5302_/A1 _4365_/Z _5015_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__or2_2
X_5888_ _6539_/A1 _5902_/A2 _5888_/B _7588_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_7627_ _7627_/D _7961_/RN _7627_/CLK _7627_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
X_4839_ _5678_/A1 _7280_/A2 _7279_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_2
XFILLER_119_473 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_5_707 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7558_ _7558_/D _7875_/RN _7881_/CLK _7558_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_119_495 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6509_ _4460_/Z _6519_/A2 _6509_/B _7880_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_20_33 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7489_ _7489_/D _7503_/CLK _7489_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_136_33 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_122_605 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_107_657 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_96_37 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_88_552 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
Xhold31 hold31/I hold31/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
Xhold20 hold20/I hold20/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
XFILLER_88_563 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_76_725 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_478 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
Xhold53 hold53/I hold53/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
Xhold64 hold64/I hold64/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
XFILLER_76_758 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_76_747 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
Xhold42 hold42/I hold42/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
XFILLER_152_76 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
Xhold86 hold86/I hold86/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
Xhold75 hold75/I hold75/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
Xhold97 hold97/I hold97/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
XFILLER_29_641 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_56_460 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_83_290 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_45_96 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XPHY_352 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_341 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_330 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_71_496 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_12_530 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_363 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_157_513 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_129_215 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_145_708 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_61_73 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_12_596 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_12_585 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_8_534 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_177_73 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_138_771 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_113_638 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_3_283 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_140_479 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_121_660 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_94_544 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_94_566 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_94_555 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_75_780 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_23_806 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6860_ _7476_/Q _6880_/C2 _6892_/A2 _7385_/Q _6860_/C _6873_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi221_1
X_6791_ _6791_/A1 _6791_/A2 _6791_/A3 _6792_/C VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_62_463 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_34_176 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5811_ _4454_/Z _5811_/A2 _5811_/B _7547_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_5742_ _5742_/A1 _5506_/C _5550_/C _5742_/A4 _5743_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor4_1
XFILLER_34_187 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5673_ _5673_/A1 _5673_/A2 _5673_/A3 _5673_/A4 _5754_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand4_1
XFILLER_175_354 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4624_ _4652_/A1 hold565/Z _4624_/B hold566/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_7412_ _7412_/D _7303_/Z _4398_/I1 _7412_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
X_7343_ _7343_/D _7298_/Z _4415_/A2 _7343_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
Xhold501 hold501/I _5922_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
X_4555_ hold781/Z _4558_/A2 _4556_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
Xhold523 _7724_/Q hold523/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
Xhold545 _7672_/Q hold545/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
XFILLER_104_605 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xhold512 hold512/I _7674_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
Xhold534 hold534/I _6496_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
Xhold567 _7951_/Q hold567/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
X_7274_ _7518_/Q _7274_/A2 _7276_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
Xhold578 _7336_/Q hold578/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
X_4486_ hold2/Z _4753_/I1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_116_487 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
Xhold556 hold556/I _7736_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
X_6225_ hold2/Z _6225_/A2 _6225_/B hold3/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
Xhold589 _7778_/Q hold589/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
X_6156_ hold302/Z _6157_/A2 hold303/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_106_69 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_850 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_861 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_5107_ _5319_/C _5692_/B _5563_/B2 _5591_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor3_2
XTAP_872 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_883 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_894 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_58_747 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_6087_ _4481_/I _6089_/A2 _6087_/B hold714/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_122_46 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_5038_ _5038_/A1 _5038_/A2 _5038_/A3 _5106_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_73_739 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_38_460 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_57_279 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_72_238 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_65_290 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_26_666 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_81_783 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_53_485 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_80_293 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_41_658 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_53_496 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6989_ _7895_/Q _7197_/A2 _6938_/I _7855_/Q _6990_/A4 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_179_693 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_166_321 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_40_179 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_31_32 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_181_357 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_135_763 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_103_2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_162_560 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_150_700 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_122_402 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_150_744 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xinput110 wb_adr_i[23] _5224_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__buf_2
Xinput154 wb_dat_i[4] _7262_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyb_1
Xinput121 wb_adr_i[4] _3728_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__buf_12
Xinput143 wb_dat_i[23] _7274_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyb_1
Xinput132 wb_dat_i[13] _7265_/B1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XFILLER_76_522 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_76_566 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_76_555 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
Xinput165 wb_stb_i _4366_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XFILLER_36_408 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_91_514 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_17_611 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_29_471 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_16_132 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_44_430 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_44_463 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_16_176 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_160 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_193 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_182 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_171 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_157_354 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_75_6 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_126_730 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_125_240 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4340_ _4340_/I _7518_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_98_124 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_87_809 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4271_ _4271_/A1 _4271_/A2 _4271_/A3 _4281_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_140_276 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_98_179 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6010_ hold583/Z _6021_/A2 _6011_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_94_374 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7961_ _7961_/D _7961_/RN _7961_/CLK _7961_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
X_6912_ _6953_/A1 _6950_/A1 _6955_/A4 _7200_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor3_4
XFILLER_47_290 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7892_ _7892_/D _7900_/RN _7892_/CLK _7892_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
X_6843_ _6843_/A1 _6843_/A2 _6843_/A3 _6848_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_63_783 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_35_496 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_149_811 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3986_ _7721_/Q hold90/I _6248_/A1 _7763_/Q _3989_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_6774_ _7720_/Q _6881_/A2 _6881_/B1 _7696_/Q _6776_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_148_321 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_5725_ _5725_/A1 _5725_/A2 _5725_/A3 _5726_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_22_179 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_5656_ _5656_/A1 _5656_/A2 _5748_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_4607_ hold866/Z _4608_/A2 _4608_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_163_357 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
Xhold320 _7989_/I hold320/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
X_5587_ _5062_/Z _5425_/B _5587_/B _5587_/C _5733_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi211_2
XFILLER_117_763 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_7326_ _7901_/RN _4334_/Z _7326_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__and2_1
X_4538_ _4460_/Z _4548_/A2 _4538_/B _7377_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
Xhold353 _7617_/Q hold353/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
Xhold331 hold331/I _7697_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
XFILLER_116_262 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xhold342 hold342/I _7609_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
XFILLER_89_113 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4469_ hold15/Z hold934/Z _4469_/B hold16/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_4
X_7257_ _7257_/A1 _7280_/A2 _7277_/B _7257_/C _7258_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi211_1
Xhold386 _7381_/Q hold386/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
XFILLER_171_390 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xhold375 _7458_/Q hold375/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
XFILLER_132_744 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_117_68 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_89_146 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_77_17 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
Xhold364 hold364/I _6075_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
Xhold397 _7730_/Q hold397/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
XFILLER_132_788 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_6208_ _6553_/A1 _6208_/A2 _6208_/B hold215/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_133_12 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7188_ _7757_/Q _7188_/A2 _7198_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_6139_ hold210/Z _6140_/A2 hold211/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_100_630 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_680 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_691 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_58_566 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_73_514 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_73_503 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_39_780 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1824 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1813 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1802 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_26_463 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_26_452 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1857 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1846 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1835 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1879 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1868 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_167_641 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_41_499 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_139_354 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_127_516 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_158_64 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_182_699 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_181_176 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
Xclkbuf_leaf_5_csclk clkbuf_leaf_9_csclk/I _7897_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_110_405 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_150_585 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_91_333 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_17_452 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_45_783 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_51_219 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_83_93 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_17_496 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_44_271 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_44_282 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3840_ _3801_/Z hold37/Z hold81/Z _3864_/A4 _4141_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand4_4
XFILLER_177_438 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3771_ hold964/Z hold966/Z _3772_/S _7967_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_158_652 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_5510_ _5621_/B _5510_/A2 _5510_/B _5752_/C _5514_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XFILLER_173_611 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6490_ _4454_/Z _6502_/A2 _6490_/B _7871_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_145_368 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_145_357 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5441_ _5591_/A2 _5501_/A2 _5613_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_66_2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_8_183 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_172_176 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5372_ _5375_/A4 _5382_/A3 _5372_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__or2_1
XFILLER_99_400 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4323_ input58/Z _4383_/A1 _4323_/B _4325_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_114_744 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7111_ _7111_/I _7115_/C VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_114_788 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_7042_ _7897_/Q _7197_/A2 _7195_/C1 _7873_/Q _7043_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_86_105 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_99_499 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4254_ _7846_/Q _6435_/A1 _4609_/A1 _7407_/Q _4256_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_4185_ _7879_/Q _6503_/A1 _6486_/A1 _7871_/Q _6124_/A1 _7701_/Q _4186_/A2 VDD VSS
+ gf180mcu_fd_sc_mcu7t5v0__aoi222_1
XFILLER_83_812 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_28_717 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_28_739 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_7944_ _7944_/D _7949_/CLK _7944_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_43_709 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1109 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_7875_ _7875_/D _7875_/RN _7875_/CLK _7875_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
X_6826_ _6826_/A1 _6767_/C _6826_/B _7433_/Q _6827_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XFILLER_51_775 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_168_449 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_149_641 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6757_ _7133_/S _6757_/A2 _6757_/B _7924_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_10_105 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_23_488 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_23_499 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_176_460 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5708_ _5104_/B _5708_/A2 _5708_/B _5710_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_3969_ _7891_/Q _6520_/A1 _5920_/A1 _7609_/Q _3981_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_6688_ _7775_/Q _6891_/C1 _6692_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_5639_ _5656_/A1 _5639_/A2 _5639_/B _5639_/C _5640_/B2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XFILLER_128_34 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_151_316 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_117_582 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xhold161 hold161/I _6460_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
Xhold150 hold150/I hold150/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
X_7309_ _7900_/RN _4334_/Z _7309_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__and2_1
Xhold183 _7378_/Q hold183/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
XFILLER_144_33 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_105_766 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
Xhold172 hold172/I _7889_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
Xhold194 hold194/I hold194/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
XFILLER_120_747 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_104_276 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_100_460 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_92_108 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_86_672 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_58_363 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2311 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2300 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_170_2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2344 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2333 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2322 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2377 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2355 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2366 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1632 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1621 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1610 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_61_539 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_27_783 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2399 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2388 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1676 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1665 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1654 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1643 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1687 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1698 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_41_274 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_174_408 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_139_140 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_167_493 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_10_672 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_127_357 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_182_474 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_154_176 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_127_379 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_6_676 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_5_164 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_5_153 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_182_496 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_154_198 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_154_187 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_142_338 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_123_574 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_68_105 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_96_458 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_77_672 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_65_812 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_37_503 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_91_141 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_80_804 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_64_366 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5990_ _6539_/A1 _6004_/A2 _5990_/B _7636_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_25_709 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4941_ _5210_/A3 _4974_/A3 _4941_/B _4941_/C _4951_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi211_4
X_7660_ _7660_/D _7877_/RN _7849_/CLK _7660_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffsnq_1
X_4872_ _4454_/Z _4872_/A2 _4872_/B hold931/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_178_747 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3823_ hold27/Z hold38/Z _6039_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_4
X_6611_ _7915_/Q _6611_/A2 _6611_/B _6612_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_165_408 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_20_458 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7591_ hold97/Z _7900_/RN _7892_/CLK hold95/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
X_3754_ _7975_/Q _7974_/Q _4291_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_2
XFILLER_158_460 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_146_600 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6542_ hold590/Z _6553_/A2 hold591/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_173_430 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_145_121 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_3685_ _7817_/Q _3685_/ZN VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_6473_ _4454_/Z _6485_/A2 _6473_/B _7863_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
Xoutput200 _4391_/ZN mgmt_gpio_oeb[36] VDD VSS gf180mcu_fd_sc_mcu7t5v0__buf_4
XFILLER_145_176 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5424_ _5424_/A1 _5575_/A2 _5424_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_173_496 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xoutput233 _8005_/Z mgmt_gpio_out[31] VDD VSS gf180mcu_fd_sc_mcu7t5v0__buf_4
Xoutput211 _7988_/Z mgmt_gpio_out[11] VDD VSS gf180mcu_fd_sc_mcu7t5v0__buf_4
XFILLER_114_530 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
Xoutput222 _7995_/Z mgmt_gpio_out[21] VDD VSS gf180mcu_fd_sc_mcu7t5v0__buf_4
Xoutput244 _7987_/Z mgmt_gpio_out[7] VDD VSS gf180mcu_fd_sc_mcu7t5v0__buf_4
X_5355_ _5680_/A1 _5768_/A3 _5546_/B1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_87_403 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
Xoutput255 _4420_/I pad_flash_io1_ie VDD VSS gf180mcu_fd_sc_mcu7t5v0__buf_4
Xoutput266 _7562_/Q pll_div[4] VDD VSS gf180mcu_fd_sc_mcu7t5v0__buf_4
Xoutput277 _7362_/Q pll_trim[15] VDD VSS gf180mcu_fd_sc_mcu7t5v0__buf_4
X_4306_ _4306_/A1 _4306_/A2 _4306_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_160_179 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5286_ _4996_/Z _5424_/A1 _5733_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_102_747 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_102_736 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_87_425 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_87_414 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
Xoutput288 _7570_/Q pll_trim[25] VDD VSS gf180mcu_fd_sc_mcu7t5v0__buf_4
Xoutput299 _4429_/Z ser_rx VDD VSS gf180mcu_fd_sc_mcu7t5v0__buf_4
XFILLER_101_224 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7025_ _7025_/A1 _7025_/A2 _7025_/A3 _7025_/A4 _7026_/A4 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand4_1
X_4237_ _7684_/Q _6090_/A1 _5874_/A1 _7585_/Q _4240_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_74_108 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_68_683 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_56_812 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xclkbuf_3_5__f_wb_clk_i clkbuf_0_wb_clk_i/Z _7959_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_114_69 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_4168_ _7613_/Q _5937_/A1 _4831_/A1 _7505_/Q _4848_/A1 _7510_/Q _4170_/A2 VDD VSS
+ gf180mcu_fd_sc_mcu7t5v0__aoi222_1
XFILLER_55_333 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4099_ _7776_/Q _6282_/A1 _6469_/A1 _7864_/Q _4100_/A4 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_7927_ _7927_/D _7938_/RN _7938_/CLK _7927_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
X_7858_ _7858_/D _7901_/RN _7858_/CLK _7858_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_70_358 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_24_742 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6809_ _7844_/Q _6894_/A2 _6891_/A2 _7828_/Q _6812_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_11_414 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_23_274 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_24_797 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7789_ _7789_/D _7901_/RN _7869_/CLK _7789_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_11_425 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_139_55 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_137_611 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_125_806 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_109_357 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xclkbuf_leaf_70_csclk _7528_/CLK _7960_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_164_463 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_152_614 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_137_699 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_136_176 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_152_658 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_2_123 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_105_596 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_105_585 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_78_425 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_2_189 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
Xclkbuf_leaf_85_csclk _7528_/CLK _7477_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_93_428 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_47_801 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_47_812 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_101_780 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_86_480 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_73_152 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_73_141 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_62_804 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_37 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_19_558 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2152 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2141 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2130 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_46_388 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_46_399 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
Xclkbuf_leaf_23_csclk _7422_/CLK _7381_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XTAP_2185 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2174 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2163 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1451 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1440 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_15_753 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_2196 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_159_224 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1484 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1473 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1462 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_30_723 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_175_706 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1495 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_175_728 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_167_290 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xclkbuf_leaf_38_csclk _7422_/CLK _7752_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_128_666 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_127_154 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
Xhold908 hold908/I _4509_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
Xhold919 _7685_/Q hold919/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
XFILLER_182_293 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_182_282 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_155_496 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_127_176 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_89_70 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_170_455 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_131_809 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_89_81 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5140_ _5543_/C _5498_/A2 _5498_/B _5187_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor3_1
XFILLER_142_179 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_97_712 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_96_211 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_69_425 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5071_ _5608_/A1 _5608_/B _5475_/B _5066_/Z _5071_/C _5072_/C VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi221_1
XFILLER_150_190 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_97_767 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_29_2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4022_ input39/Z _5903_/A1 _6316_/A1 _7794_/Q _4024_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_38_812 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_56_108 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5973_ hold47/Z _5987_/A2 _5973_/B _7628_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_92_494 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4924_ _4924_/A1 _4924_/A2 _4924_/A3 _4924_/A4 _4926_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand4_1
X_7712_ _7712_/D _7853_/RN _7812_/CLK _7712_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_178_522 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_21_712 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7643_ _7643_/D _7923_/RN _7792_/CLK _7643_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
X_4855_ hold47/Z _4857_/A2 _4855_/B hold414/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_159_780 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3806_ _3810_/S hold148/Z _3806_/B _3864_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi21_4
XFILLER_119_622 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_119_611 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7574_ hold23/Z _7875_/RN _7847_/CLK _7982_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
X_4786_ _7219_/A1 _4795_/S _4786_/B _7478_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_181_709 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3737_ _7346_/Q _7344_/Q _3774_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_119_633 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_118_132 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_6525_ hold593/Z _6536_/A2 hold594/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_146_463 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_107_806 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3668_ _7951_/Q _7248_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_173_293 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_161_411 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_133_124 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_133_102 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_118_176 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6456_ _4454_/Z _6468_/A2 _6456_/B _7855_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_5407_ _5782_/A1 _5407_/A2 _5407_/A3 _5414_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand3_1
X_6387_ hold896/Z _6400_/A2 _6388_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_161_499 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5338_ _5338_/A1 _5421_/B1 _5779_/B1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_125_35 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_649 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7008_ _7008_/A1 _7008_/A2 _7008_/A3 _7008_/A4 _7026_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand4_1
X_5269_ _5624_/A1 _5624_/B _5586_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_75_428 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_29_812 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_71_601 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_28_388 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_141_89 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_169_511 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_169_566 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_70_188 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_157_728 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_133_2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_7_215 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_165_783 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_152_400 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_137_485 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_125_636 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_180_764 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_113_809 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_124_179 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_79_712 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_509 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_3_487 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_79_767 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_59_73 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_78_277 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_38_108 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_115_90 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_47_686 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_179_319 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_61_144 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_15_550 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1292 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1281 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1270 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_30_531 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_147_227 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4640_ _4652_/A1 _4640_/A2 _4640_/B hold485/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_175_558 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_163_709 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_128_463 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6310_ hold725/Z _6315_/A2 _6311_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_4571_ _6539_/A1 _4573_/A2 _4571_/B _7391_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_143_422 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_143_411 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_143_400 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7290_ _7901_/RN _4334_/Z _7290_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__and2_1
Xhold727 _7835_/Q hold727/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
Xhold705 _7690_/Q hold705/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
Xhold716 _7353_/Q hold716/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
XFILLER_171_753 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6241_ _7755_/Q hold6/Z _6242_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_143_444 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_143_455 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xhold738 _7476_/Q hold738/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
Xhold749 _7546_/Q hold749/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
X_6172_ _4481_/I _6174_/A2 _6172_/B _7722_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_143_499 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_130_105 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5123_ _4953_/Z _5139_/A1 _5014_/Z _5543_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand3_4
X_5054_ _5199_/B _3727_/I _5054_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__or2_2
XFILLER_69_288 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_57_428 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_84_258 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4005_ _7882_/Q _6503_/A1 _6005_/A1 _7648_/Q _4024_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_37_141 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_93_792 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_53_601 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_25_347 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_5956_ hold47/Z _5970_/A2 _5956_/B _7620_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_178_352 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4907_ _5302_/A1 _5224_/A3 _5224_/A4 _5016_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor3_4
X_5887_ hold740/Z _5902_/A2 _5888_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_52_188 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4838_ _7516_/Q _5301_/B _5520_/C VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_4
X_7626_ _7626_/D _7961_/RN _7960_/CLK _7626_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_119_463 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4769_ _4769_/A1 _6537_/A2 _4773_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_7557_ _7557_/D _7875_/RN _7563_/CLK _7557_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffsnq_1
XFILLER_147_783 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_146_282 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6508_ hold677/Z _6519_/A2 _6509_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_7488_ _7488_/D _7503_/CLK _7488_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_6439_ _4454_/Z _6451_/A2 _6439_/B _7847_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_121_116 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_121_105 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_106_179 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_161_296 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_115_691 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_88_531 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xhold10 hold10/I hold10/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
Xhold32 hold32/I hold32/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
Xhold21 hold21/I hold21/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
XFILLER_0_457 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xhold54 hold54/I hold54/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
Xhold43 hold43/I hold43/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
Xhold65 hold65/I hold65/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
Xhold87 hold87/I hold87/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
Xhold98 hold98/I hold98/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
Xhold76 hold76/I hold76/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
XFILLER_29_98 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_43_144 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_45_86 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_342 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_331 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_320 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_364 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_353 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_12_575 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_8_524 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_125_499 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_112_105 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_112_116 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_121_650 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_67_704 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_94_534 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_39_428 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_120_193 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_66_247 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_19_141 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_81_228 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_19_152 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_34_133 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_47_494 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6790_ _7753_/Q _6644_/Z _6885_/B1 _7713_/Q _6791_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_5810_ hold867/Z _5811_/A2 _5811_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_5741_ _5741_/A1 _4993_/B _5741_/A3 _5741_/B _5742_/A4 VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai31_1
XFILLER_96_2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_22_339 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_34_199 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_176_812 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7411_ _7411_/D _7302_/Z _4415_/A2 _7411_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffsnq_2
X_5672_ _5179_/B _5672_/A2 _5793_/A2 _5606_/B _5673_/A4 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_4623_ hold564/Z _3830_/Z _4623_/B hold565/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_7342_ _7342_/D _7297_/Z _4415_/A2 _7342_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_129_783 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xhold502 hold502/I _7604_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
X_4554_ _4554_/A1 _6537_/A2 _4558_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_7273_ _7273_/A1 _7277_/B _7273_/B _7956_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_144_742 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
Xhold524 _7720_/Q hold524/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
Xhold513 _7620_/Q hold513/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
Xhold535 hold535/I _7874_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
X_4485_ hold1/Z hold934/Z _4485_/B hold935/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_4
Xhold557 _7460_/Q hold557/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
Xhold568 hold568/I _4627_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
X_6224_ _7747_/Q _6225_/A2 _6225_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
Xhold579 _3793_/Z hold579/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
XFILLER_116_477 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xhold546 hold546/I _6066_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
XFILLER_131_425 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_103_138 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6155_ _4481_/I _6157_/A2 _6155_/B hold663/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_106_59 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_106_37 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_100_812 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_840 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_851 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_862 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_5106_ _5106_/A1 _5106_/A2 _5106_/A3 _5106_/A4 _5115_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor4_1
X_6086_ hold712/Z _6089_/A2 hold713/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_873 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_884 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_895 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_5037_ _5585_/A1 _5658_/B _5608_/B _5669_/A1 _5037_/C _5038_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi221_1
XFILLER_85_567 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_73_729 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_66_792 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_26_612 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_80_250 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_25_155 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_25_144 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_26_689 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6988_ _7887_/Q _7196_/A2 _7196_/B1 _7637_/Q _6990_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_167_812 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_139_503 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5939_ hold47/Z _5953_/A2 _5939_/B _7612_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_166_377 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_7609_ _7609_/D _7923_/RN _7792_/CLK _7609_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_21_394 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_135_753 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_1_700 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_163_21 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_150_756 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_107_499 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xinput100 wb_adr_i[14] _4922_/A4 VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyc_1
Xinput111 wb_adr_i[24] _4370_/A4 VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XFILLER_163_54 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_122_458 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
Xinput144 wb_dat_i[24] _7240_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyb_1
Xinput133 wb_dat_i[14] _7269_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyb_1
Xinput122 wb_adr_i[5] _5369_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__buf_12
XFILLER_130_480 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_102_160 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_76_534 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
Xinput166 wb_we_i _3658_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
Xinput155 wb_dat_i[5] _7267_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XFILLER_0_298 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_48_247 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_63_228 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_56_63 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_17_634 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_112_91 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_71_283 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_176_108 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_158_812 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_161 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_150 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_9_800 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XPHY_194 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_183 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_172 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_8_321 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_145_517 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_12_383 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_8_343 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_157_388 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_126_720 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_141_712 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_113_425 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_4_593 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4270_ _7870_/Q _6486_/A1 _5849_/A2 _7572_/Q _4271_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_95_810 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_100_108 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_67_567 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_11_2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7960_ _7960_/D _7961_/RN _7960_/CLK _7960_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_48_770 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7891_ _7891_/D _7901_/RN _7896_/CLK _7891_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
X_6911_ _6599_/Z _6941_/A2 _6908_/Z _7191_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor3_4
X_6842_ _7765_/Q _6892_/A2 _6892_/B1 _7731_/Q _6843_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_62_250 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_22_114 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_23_637 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_23_626 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3985_ _3985_/A1 _3985_/A2 _3985_/A3 _3985_/A4 _3990_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand4_1
X_6773_ _7656_/Q _6882_/B1 _6647_/Z _7616_/Q _6776_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_5724_ _5759_/A1 _5724_/A2 _5724_/B _5725_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_176_664 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_175_130 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_175_141 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5655_ _5766_/A1 _5804_/A1 _5655_/A3 _5655_/A4 _5676_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor4_1
XFILLER_109_709 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4606_ _6539_/A1 _4608_/A2 _4606_/B _7405_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_7325_ _7877_/RN _4334_/Z _7325_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__and2_1
Xhold310 hold310/I _6502_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
X_5586_ _5586_/A1 _5586_/A2 _5586_/A3 _5586_/A4 _5589_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand4_1
X_4537_ hold689/Z _4548_/A2 _4538_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
Xhold321 hold321/I _4706_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
Xhold332 _7689_/Q hold332/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
Xhold343 _7803_/Q hold343/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
Xhold387 _7952_/Q hold387/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
X_7256_ _7256_/A1 _7256_/A2 _7257_/C VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_4468_ hold49/I _7263_/A1 _4469_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
Xhold376 hold376/I _4744_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
XFILLER_132_734 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
Xhold354 hold354/I _7617_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
XFILLER_117_47 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xhold365 hold365/I _7676_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
X_6207_ hold213/Z _6208_/A2 hold214/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
Xhold398 _7527_/Q hold398/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
X_7187_ _7133_/S _7187_/A2 _7187_/B _7939_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_4399_ _7436_/Q input67/Z _7335_/Q _4399_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_6138_ _4481_/I _6140_/A2 _6138_/B hold499/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
XTAP_670 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_58_501 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_58_534 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_133_46 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_681 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_692 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_133_68 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_93_17 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6069_ hold510/Z _6072_/A2 hold511/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_39_792 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_54_740 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1825 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1814 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1803 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_54_751 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1858 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1847 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1836 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_81_570 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_26_486 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_53_283 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_158_108 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1869 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_13_158 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_41_445 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_41_456 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_13_169 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_10_810 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_22_670 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_167_664 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_166_141 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_158_32 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_158_76 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_182_667 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_181_144 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_135_550 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_123_712 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_107_241 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_5_357 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_150_531 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_123_778 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_96_629 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_122_277 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_95_139 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_67_73 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_37_707 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_49_567 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_44_250 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_83_83 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_177_428 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_32_434 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3770_ hold965/Z hold62/I _3772_/S _7968_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_157_141 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_157_130 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_9_641 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5440_ _5705_/B _5712_/B _5555_/B _5534_/A2 _5444_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor4_1
XFILLER_8_195 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5371_ _5371_/A1 _5371_/A2 _5371_/B _5371_/C _5382_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_59_2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4322_ _4322_/A1 _4322_/A2 _7337_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_126_594 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_7110_ _7714_/Q _7189_/A2 _7191_/B1 _7804_/Q _7111_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_7041_ _7833_/Q _7203_/A2 _6938_/I _7857_/Q _7043_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_99_456 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4253_ _4253_/A1 _4253_/A2 _4253_/A3 _4253_/A4 _4263_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand4_1
XFILLER_141_586 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_101_428 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4184_ input47/Z _4231_/B1 _5817_/A1 _7559_/Q _5807_/A1 _7547_/Q _4186_/A1 VDD VSS
+ gf180mcu_fd_sc_mcu7t5v0__aoi222_1
Xclkbuf_3_4__f_wb_clk_i clkbuf_0_wb_clk_i/Z _7545_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_55_515 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_94_183 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_82_312 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_7943_ _7943_/D _7949_/CLK _7943_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_82_389 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_63_570 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7874_ _7874_/D _7875_/RN _7874_/CLK _7874_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_35_283 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6825_ _6825_/A1 _6825_/A2 _6825_/A3 _6826_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor3_1
XFILLER_35_294 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3968_ _7827_/Q _6384_/A1 _3968_/B _3981_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_6756_ _7924_/Q _7133_/S _6757_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_51_798 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5707_ _5782_/A2 _5704_/Z _5706_/Z _5717_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand3_1
X_3899_ _7789_/Q _6299_/A1 _6435_/A1 _7853_/Q _3901_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_6687_ _7799_/Q _6883_/A2 _6883_/B1 _7783_/Q _6705_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_163_144 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5638_ _5064_/B _5678_/A3 _5637_/Z _7279_/B _5639_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai31_1
XFILLER_163_177 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5569_ _5376_/B _5218_/C _5587_/C VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_105_712 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_88_17 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_88_28 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xhold162 hold162/I _7857_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
Xhold151 hold151/I _7566_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
Xhold140 hold140/I _7627_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
X_7308_ _7875_/RN _4334_/Z _7308_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__and2_1
Xhold184 _7683_/Q hold184/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
Xhold173 _7761_/Q hold173/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
XFILLER_105_778 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
Xhold195 hold195/I _7350_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
X_7239_ _7518_/Q _7239_/A2 _7241_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_144_56 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_132_575 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_104_266 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_85_161 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_85_150 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_18_206 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2301 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_73_312 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2334 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2323 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2312 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1600 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_61_507 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_37_98 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2378 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2356 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2367 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2345 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_163_2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1633 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1622 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1611 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_26_250 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_2389 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1666 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1655 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1644 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_159_428 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1688 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1699 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1677 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_41_264 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_41_286 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_96_404 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_110_203 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_111_759 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_110_247 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_110_269 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_92_676 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_52_507 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_52_518 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4940_ _4946_/A1 _5230_/A1 _5200_/B _4974_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_4
XFILLER_91_164 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_64_389 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_18_784 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_45_570 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_52_529 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_17_283 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4871_ hold929/Z _4872_/A2 hold930/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_33_732 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_3822_ _3801_/Z hold37/Z _3843_/A3 _3864_/A4 hold38/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand4_4
X_7590_ _7590_/D _7900_/RN _7592_/CLK _8000_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
X_6610_ _7434_/Q _7915_/Q _6610_/A3 _6611_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_177_247 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_20_448 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6541_ _4454_/Z _6553_/A2 _6541_/B _7895_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_3753_ _4383_/A1 _7413_/Q _4292_/B _3772_/S VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand3_4
X_3684_ _7825_/Q _3684_/ZN VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_118_347 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6472_ hold874/Z _6485_/A2 _6473_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
Xoutput201 _4389_/ZN mgmt_gpio_oeb[37] VDD VSS gf180mcu_fd_sc_mcu7t5v0__buf_4
XFILLER_145_144 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5423_ _5624_/A1 _5648_/B2 _5724_/B _5627_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
Xoutput234 _4394_/Z mgmt_gpio_out[32] VDD VSS gf180mcu_fd_sc_mcu7t5v0__buf_4
X_5354_ _5354_/A1 _5354_/A2 _5354_/A3 _5354_/A4 _5356_/A4 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor4_1
Xoutput212 _7989_/Z mgmt_gpio_out[12] VDD VSS gf180mcu_fd_sc_mcu7t5v0__buf_4
Xoutput223 _7996_/Z mgmt_gpio_out[22] VDD VSS gf180mcu_fd_sc_mcu7t5v0__buf_4
X_4305_ _7414_/Q _4308_/S _7340_/Q _4306_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
Xoutput245 _4399_/Z mgmt_gpio_out[8] VDD VSS gf180mcu_fd_sc_mcu7t5v0__buf_4
Xoutput267 _7556_/Q pll_ena VDD VSS gf180mcu_fd_sc_mcu7t5v0__buf_4
Xoutput256 _4420_/ZN pad_flash_io1_oe VDD VSS gf180mcu_fd_sc_mcu7t5v0__buf_4
X_5285_ _5663_/A1 _5692_/B _5285_/A3 _5287_/C VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor3_1
XFILLER_99_286 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_87_437 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
Xoutput289 _7365_/Q pll_trim[2] VDD VSS gf180mcu_fd_sc_mcu7t5v0__buf_4
Xoutput278 _7347_/Q pll_trim[16] VDD VSS gf180mcu_fd_sc_mcu7t5v0__buf_4
X_7024_ _7816_/Q _7207_/A2 _7207_/B1 _7718_/Q _7024_/C _7025_/A4 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi221_1
XFILLER_87_459 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4236_ _4236_/A1 _4236_/A2 _4236_/A3 _4236_/A4 _4283_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand4_2
XFILLER_114_37 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_68_673 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4167_ _4167_/A1 _4167_/A2 _4167_/A3 _4167_/A4 _4167_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__and4_1
XFILLER_82_120 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_28_526 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4098_ _7750_/Q _6226_/A1 _6401_/A1 _7832_/Q _4100_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_82_131 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_71_805 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_28_559 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7926_ _7926_/D _7938_/RN _7935_/CLK _7926_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_24_721 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_43_518 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_55_389 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_169_726 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7857_ _7857_/D _7901_/RN _7899_/CLK _7857_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
Xclkbuf_leaf_4_csclk clkbuf_leaf_9_csclk/I _7592_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
X_6808_ _7730_/Q _6892_/B1 _6880_/B1 _7812_/Q _6815_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_168_247 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7788_ _7788_/D _7900_/RN _7898_/CLK _7788_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_23_286 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_135_6 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6739_ hold78/I _6880_/C2 _6881_/B1 _7695_/Q _7809_/Q _6880_/B1 _6742_/A1 VDD VSS
+ gf180mcu_fd_sc_mcu7t5v0__aoi222_1
XFILLER_99_27 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_136_166 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_136_155 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_151_125 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_151_103 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_2_113 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_151_158 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_2_179 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_120_534 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_59_651 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_48_53 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_74_676 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_27 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_46_356 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2153 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2142 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2131 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2120 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_64_63 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_64_52 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_27_570 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2186 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2175 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2164 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1441 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1430 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_61_359 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2197 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1474 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1452 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1463 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_159_247 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1496 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1485 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_80_51 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_30_735 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_127_166 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_127_144 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
Xhold909 hold909/I _7364_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
XFILLER_6_463 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_170_445 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_89_93 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_123_350 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_69_404 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5070_ _5458_/C _5527_/A1 _5458_/B _5071_/C VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor3_1
XFILLER_111_534 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_111_567 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_97_779 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4021_ _7866_/Q _6469_/A1 _6418_/A1 _7842_/Q _4024_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_49_150 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_77_481 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_37_312 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_53_805 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_5972_ hold490/Z _5987_/A2 _5973_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_80_624 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_80_602 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4923_ _4923_/A1 input97/Z _4926_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_7711_ hold86/Z _7853_/RN _7722_/CLK hold84/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_178_534 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_60_392 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4854_ hold412/Z _4857_/A2 hold413/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_7642_ _7642_/D _7961_/RN _7961_/CLK _7642_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
X_3805_ hold36/Z _3803_/Z _3810_/S hold37/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_7573_ _7573_/D _7901_/RN _7829_/CLK _7573_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_20_245 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_21_779 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4785_ _7478_/Q _4795_/S _4786_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_3736_ _7976_/Q _3734_/Z _3736_/B _3741_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_118_122 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6524_ _4454_/Z _6536_/A2 _6524_/B _7887_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_118_166 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_173_283 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3667_ hold45/I _7243_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_161_423 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6455_ hold879/Z _6468_/A2 _6456_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_161_445 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5406_ _5292_/B _5779_/B1 _5587_/B _5406_/C _5407_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi211_1
X_6386_ _6539_/A1 _6400_/A2 _6386_/B _7822_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_5337_ _5680_/A1 _5779_/A2 _5680_/B1 _5680_/B2 _5337_/C _5343_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi221_1
XFILLER_87_212 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_142_692 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_125_47 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5268_ _5394_/A1 _5005_/Z _5687_/B _5645_/A3 _5680_/C VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor4_2
XFILLER_102_534 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_102_567 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_87_278 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_7007_ _7710_/Q _7189_/A2 _7191_/B1 _7800_/Q _7008_/A4 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_4219_ input11/Z _4219_/A2 _5812_/A1 _7556_/Q _4262_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_5199_ _4915_/Z _4996_/Z _5199_/B _5371_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_18_34 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_141_46 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_56_654 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_16_529 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_56_676 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_71_668 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_70_112 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7909_ _7909_/D _7938_/RN _7940_/CLK _7909_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_4
XFILLER_24_540 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_12_724 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_11_212 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_34_66 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_8_717 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_126_2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_164_250 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_109_144 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_166_76 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_164_272 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_109_177 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_166_98 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_121_810 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_112_309 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_133_692 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_79_757 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_3_499 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_78_256 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_93_215 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_59_492 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_75_73 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_62_624 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_62_602 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_74_495 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_62_635 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_15_540 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1293 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1282 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1271 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1260 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_392 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4570_ hold780/Z _4573_/A2 _4571_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_155_283 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xhold717 _7867_/Q hold717/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
Xhold728 _7891_/Q hold728/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
Xhold706 hold706/I _6104_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
XFILLER_7_783 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6240_ hold233/Z hold6/Z _6240_/B hold234/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
Xhold739 _7470_/Q hold739/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
XFILLER_171_798 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_6171_ hold657/Z _6174_/A2 _6172_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_41_2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5122_ _4953_/Z _5139_/A1 _5014_/Z _5122_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__and3_1
XFILLER_97_532 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_69_212 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5053_ _5199_/B _3727_/I _5303_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_4
X_4004_ _7890_/Q _6520_/A1 _4032_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_65_451 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_1_70 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_25_304 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_38_676 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5955_ hold513/Z _5970_/A2 _5956_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_40_307 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_53_668 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4906_ _4905_/Z _5302_/A3 _4906_/S _4906_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_80_487 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5886_ _5886_/A1 _6537_/A2 _5902_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_4
XFILLER_33_370 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_40_318 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4837_ _7519_/Q _7518_/Q _7520_/Q _5301_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__or3_1
XFILLER_166_526 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xclkbuf_leaf_84_csclk _7528_/CLK _7637_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
X_7625_ _7625_/D _7961_/RN _7876_/CLK _7625_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_146_250 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4768_ _4454_/Z _4768_/A2 _4768_/B _7471_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_5_709 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7556_ _7556_/D input75/Z _7563_/CLK _7556_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_146_272 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4699_ hold476/Z _4718_/A1 hold477/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_112_8 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7487_ _7487_/D _7503_/CLK _7487_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_3719_ _7906_/Q _6633_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_3
X_6507_ _4454_/Z _6519_/A2 _6507_/B _7879_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_161_242 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6438_ hold880/Z _6451_/A2 _6439_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_136_68 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_96_17 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_403 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_161_286 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6369_ hold47/Z _6383_/A2 _6369_/B _7814_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
Xhold11 hold11/I hold11/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
XFILLER_130_673 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xhold22 hold22/I hold22/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
Xhold33 hold33/I hold33/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
XFILLER_152_34 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xhold44 hold44/I hold44/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
XFILLER_130_695 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xhold55 hold55/I hold55/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
XFILLER_76_749 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_75_215 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
Xhold66 hold66/I hold66/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
Xhold88 hold88/I hold88/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
Xhold99 hold99/I hold99/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
Xhold77 hold77/I hold77/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
Xclkbuf_leaf_37_csclk clkbuf_3_7__f_csclk/Z _7729_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_29_698 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_44_602 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_56_473 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_83_292 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_310 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_343 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_332 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_321 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
Xclkbuf_0_mgmt_gpio_in[4] mgmt_gpio_in[4] clkbuf_0_mgmt_gpio_in[4]/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XPHY_365 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_354 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_24_392 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_157_559 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_8_536 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_165_570 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_6_37 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_180_551 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_99_808 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_4_742 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_98_318 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_3_241 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_112_139 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_112_128 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_120_172 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_19_164 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_35_602 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_47_462 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_22_307 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_50_605 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5740_ _5740_/A1 _5740_/A2 _5740_/A3 _5739_/Z _5804_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand4_1
XFILLER_15_381 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_22_318 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1090 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_5671_ _5774_/C _5671_/A2 _5748_/A2 _5671_/A4 _5671_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__or4_1
XFILLER_89_2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7410_ _7410_/D _7875_/RN _7410_/CLK _7410_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
X_4622_ _3830_/Z hold47/Z _4623_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_7341_ _7341_/D _7296_/Z _4415_/A2 _7341_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_128_250 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4553_ _4454_/Z _4553_/A2 _4553_/B _7384_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_7272_ _7272_/A1 _7280_/A2 _7277_/B _7272_/C _7273_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi211_1
X_4484_ hold49/I _7278_/A1 _4485_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_171_540 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
Xhold514 _7424_/Q hold514/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
XFILLER_144_732 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
Xhold525 _7696_/Q hold525/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
Xhold536 _7688_/Q hold536/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
Xhold503 _7738_/Q hold503/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
Xhold569 hold569/I hold569/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
X_6223_ hold233/Z _6225_/A2 _6223_/B _7746_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
Xhold558 hold558/I hold558/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
XFILLER_143_242 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xhold547 hold547/I _7672_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
XFILLER_143_286 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6154_ hold661/Z _6157_/A2 hold662/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_830 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_841 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_852 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_6085_ _4476_/I _6089_/A2 _6085_/B hold347/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_112_673 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5105_ _5105_/A1 _5105_/A2 _5105_/A3 _5105_/A4 _5106_/A4 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand4_1
XFILLER_85_524 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_863 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_874 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_885 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_57_215 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5036_ _5714_/A1 _5797_/A1 _5099_/B _5037_/C VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XTAP_896 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_122_37 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_26_602 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6987_ _7645_/Q _7195_/A2 _7195_/B1 _7621_/Q _7195_/C1 _7871_/Q _6990_/A2 VDD VSS
+ gf180mcu_fd_sc_mcu7t5v0__aoi222_1
XFILLER_53_443 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_53_465 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_53_454 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_15_35 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5938_ hold670/Z _5953_/A2 _5939_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_40_115 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_41_638 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_80_295 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_178_194 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5869_ _7581_/Q _5870_/A1 _5870_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_154_507 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7608_ _7608_/D _7923_/RN _7736_/CLK _7608_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_166_389 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_147_570 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_147_12 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7539_ _7539_/D _7959_/RN _7545_/CLK hold70/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_107_412 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_119_283 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_31_89 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_162_551 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_122_415 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_1_712 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xinput101 wb_adr_i[15] _4922_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyc_1
XFILLER_0_244 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xinput145 wb_dat_i[25] _7245_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyb_1
Xinput134 wb_dat_i[15] _7275_/B1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyb_1
Xinput112 wb_adr_i[25] _3660_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyb_1
Xinput123 wb_adr_i[6] _5199_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__buf_12
Xinput156 wb_dat_i[6] _7272_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XFILLER_76_546 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_48_237 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_72_763 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_32_605 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_151 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_140 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
Xclkbuf_3_1__f_csclk clkbuf_0_csclk/Z clkbuf_leaf_9_csclk/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_169_172 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_184 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_173 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_162 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_9_812 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_195 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_75_8 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_8_333 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_157_378 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_8_388 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_153_540 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_153_551 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_180_392 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_141_735 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_125_286 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_113_437 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_99_638 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_98_148 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_97_93 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_39_215 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
Xclkbuf_3_3__f_wb_clk_i clkbuf_0_wb_clk_i/Z _7938_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_94_321 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_55_708 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6910_ _6599_/Z _6950_/A2 _6955_/A4 _7203_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor3_4
X_7890_ _7890_/D _7900_/RN _7898_/CLK _7890_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
X_6841_ _7829_/Q _6891_/A2 _6891_/B1 _7675_/Q _6891_/C1 _7781_/Q _6843_/A2 VDD VSS
+ gf180mcu_fd_sc_mcu7t5v0__aoi222_1
XFILLER_90_560 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_50_402 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_3984_ _7713_/Q _6141_/A1 _6316_/A1 _7795_/Q _3985_/A4 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_6772_ _7648_/Q _6880_/C2 _6892_/A2 _7762_/Q _6776_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_5723_ _5723_/A1 _5723_/A2 _5791_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_50_479 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_176_676 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5654_ _5740_/A3 _5651_/Z _5654_/A3 _5655_/A4 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_175_175 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_148_389 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_129_570 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4605_ hold778/Z _4608_/A2 _4606_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_7324_ _7877_/RN _4334_/Z _7324_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_163_359 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xhold311 hold311/I _7877_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
X_5585_ _5585_/A1 _5658_/B _5585_/B _5585_/C _5586_/A4 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi211_1
Xhold300 hold300/I _6483_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
X_4536_ _4454_/Z _4548_/A2 _4536_/B _7376_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
Xhold322 hold322/I _7440_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
Xhold344 hold344/I _7803_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
Xhold333 hold333/I _6102_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
X_7255_ _7520_/Q _7255_/A2 _7255_/B1 _7519_/Q _7256_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_1
Xhold366 _7633_/Q hold366/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
Xhold377 hold377/I _7458_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
XFILLER_144_584 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_131_212 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_116_275 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
Xhold355 _7657_/Q hold355/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
XFILLER_89_126 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4467_ _4487_/A1 _6545_/A1 _4467_/B hold195/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_4398_ _7437_/Q _4398_/I1 _7334_/Q _4398_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_6206_ _4481_/I _6208_/A2 _6206_/B hold505/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
Xhold388 hold388/I _7577_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
Xhold399 hold399/I _4870_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
X_7186_ _7939_/Q _7133_/S _7187_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_6137_ hold497/Z _6140_/A2 hold498/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_660 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_671 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_682 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_693 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_58_546 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_133_58 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6068_ _4476_/I _6072_/A2 _6068_/B hold328/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_100_676 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_85_354 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_39_771 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5019_ _5200_/B _5230_/A1 _5024_/A2 _5201_/B _5021_/B1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai31_2
XFILLER_73_538 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1815 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1804 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_14_605 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_26_34 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1848 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1837 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1826 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_26_67 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1859 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_13_148 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_139_301 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_42_33 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_166_120 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_181_101 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_174_21 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_135_540 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_162_392 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_107_286 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_150_543 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_3_27 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_76_321 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_91_335 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_57_590 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_91_357 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_29_292 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_45_763 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_83_73 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_60_744 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_60_788 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_13_682 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_158_676 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_161_808 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_66_4 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5370_ _5369_/B _5381_/A2 _5370_/B _5375_/A4 VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_2
XFILLER_160_318 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4321_ _4383_/A1 _7411_/Q _7337_/Q _4322_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_114_724 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_113_212 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7040_ _7825_/Q _7202_/A2 _7201_/B1 _7671_/Q _7043_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_4_380 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4252_ _7387_/Q _4559_/A1 _4779_/A1 _7476_/Q _4253_/A4 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_95_641 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4183_ _4183_/A1 _4183_/A2 _4183_/A3 _4187_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_94_151 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_103_17 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7942_ _7942_/D _7949_/CLK _7942_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_27_229 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7873_ _7873_/D _7901_/RN _7873_/CLK _7873_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_23_413 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6824_ _6824_/A1 _6824_/A2 _6824_/A3 _6824_/A4 _6825_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand4_1
XFILLER_168_429 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_3967_ _4075_/B _4155_/A2 _3968_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_6755_ _7433_/Q _7923_/Q _6755_/B _6757_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_5706_ _5706_/A1 _5706_/A2 _5706_/A3 _5706_/A4 _5706_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__and4_1
XFILLER_164_602 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3898_ _7611_/Q _5920_/A1 _5971_/A1 _7635_/Q _3901_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_6686_ _7002_/B _6686_/A2 _6686_/A3 _6686_/B _7921_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai31_1
XFILLER_148_197 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5637_ _5637_/A1 _5679_/A1 _5637_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_136_337 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_151_307 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5568_ _5104_/B _5708_/A2 _5578_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_132_521 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
Xhold130 hold130/I _7735_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
XFILLER_104_201 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4519_ hold233/Z _4521_/A2 _4519_/B hold475/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
Xhold152 _7607_/Q hold152/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
Xhold141 _7447_/Q hold141/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
X_7307_ _7875_/RN _4334_/Z _7307_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__and2_1
X_5499_ _5499_/A1 _5499_/A2 _5653_/A1 _5499_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__or3_1
X_7238_ _7279_/B _7238_/A2 _7238_/A3 _7280_/A3 _7277_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand4_4
Xhold163 _7849_/Q hold163/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
XFILLER_144_392 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xhold185 hold185/I _6089_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
Xhold174 hold174/I _6256_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
XFILLER_105_757 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xhold196 _7675_/Q hold196/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
XFILLER_86_630 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7169_ _7535_/Q _7197_/A2 _7196_/A2 _7546_/Q _7196_/B1 _7474_/Q _7172_/A1 VDD VSS
+ gf180mcu_fd_sc_mcu7t5v0__aoi222_1
XFILLER_58_321 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_490 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_37_33 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2302 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_160_34 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_100_495 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_46_538 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_58_387 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_58_398 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2335 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2324 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2313 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_160_56 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_73_357 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2357 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2368 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2346 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1623 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1612 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1601 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_14_402 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_2379 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_156_2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1667 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1656 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1645 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1634 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_744 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1689 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1678 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_139_120 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_167_451 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_154_112 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_154_123 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_182_454 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_170_605 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_143_808 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_5_144 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_142_318 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_150_351 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_111_716 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_78_62 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_77_641 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_110_259 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_77_674 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_37_516 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_49_354 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_49_376 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_49_398 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_91_121 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_64_368 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_91_176 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_33_700 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_17_295 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_4870_ hold47/Z _4872_/A2 _4870_/B hold400/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_178_749 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_177_215 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3821_ hold609/Z hold76/Z _6486_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_4
XFILLER_60_552 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_32_243 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_32_276 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_6540_ hold804/Z _6553_/A2 _6541_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_3752_ _3752_/I _3756_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_146_602 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_71_2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_146_646 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_118_337 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3683_ _7833_/Q _3683_/ZN VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_6471_ _6539_/A1 _6485_/A2 _6471_/B _7862_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_9_494 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5422_ _5660_/A2 _5422_/A2 _5422_/B _5439_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
Xoutput235 _4395_/Z mgmt_gpio_out[33] VDD VSS gf180mcu_fd_sc_mcu7t5v0__buf_4
XFILLER_161_627 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
Xoutput213 _4412_/Z mgmt_gpio_out[13] VDD VSS gf180mcu_fd_sc_mcu7t5v0__buf_4
X_5353_ _5353_/A1 _5642_/A2 _5493_/B _5353_/A4 _5354_/A4 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand4_1
Xoutput224 _7997_/Z mgmt_gpio_out[23] VDD VSS gf180mcu_fd_sc_mcu7t5v0__buf_4
Xoutput202 _3709_/ZN mgmt_gpio_oeb[3] VDD VSS gf180mcu_fd_sc_mcu7t5v0__buf_4
X_4304_ _4304_/I0 _7342_/Q _4309_/S _7342_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_126_392 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xoutput246 _4398_/Z mgmt_gpio_out[9] VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_1
Xoutput257 _7566_/Q pll90_sel[0] VDD VSS gf180mcu_fd_sc_mcu7t5v0__buf_4
Xoutput268 _7563_/Q pll_sel[0] VDD VSS gf180mcu_fd_sc_mcu7t5v0__buf_4
X_5284_ _5573_/A1 _5292_/B _5247_/B _5431_/B _5288_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_1
Xoutput279 _7348_/Q pll_trim[17] VDD VSS gf180mcu_fd_sc_mcu7t5v0__buf_4
XFILLER_101_215 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_7023_ _7023_/A1 _7023_/A2 _7023_/A3 _7024_/C VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand3_1
X_4235_ _7822_/Q _6384_/A1 _4863_/A1 _7525_/Q _4236_/A4 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_95_460 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_83_600 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_68_663 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4166_ _7364_/Q _4505_/A1 _6005_/A1 _7645_/Q _4167_/A4 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_68_685 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4097_ _7654_/Q _6022_/A1 _6537_/A1 _7896_/Q _4100_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_55_357 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_130_26 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7925_ _7925_/D _7938_/RN _7935_/CLK _7925_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_82_176 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_130_37 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7856_ _7856_/D _7901_/RN _7866_/CLK _7856_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffsnq_1
XFILLER_82_198 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_24_744 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6807_ _7796_/Q _6893_/A2 _6890_/B1 _7852_/Q _6815_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_23_254 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_51_574 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7787_ _7787_/D _7901_/RN _7833_/CLK _7787_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
X_4999_ _4999_/A1 _4999_/A2 _4999_/A3 _4999_/A4 _4999_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__and4_1
XFILLER_23_35 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6738_ _6738_/A1 _6738_/A2 _6738_/A3 _6738_/A4 _6753_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand4_1
XFILLER_23_79 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_136_112 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_128_6 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6669_ _7822_/Q _6891_/A2 _6894_/C1 _7830_/Q _6683_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_152_605 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_124_318 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_3_637 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_151_137 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_78_449 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_59_641 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_48_32 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_171_33 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_86_460 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2110 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_58_195 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2143 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2132 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2121 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2176 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2165 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2154 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1442 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1431 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1420 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2198 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2187 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_159_215 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1475 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1453 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1464 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1497 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1486 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_30_747 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_155_443 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_127_134 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_155_487 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_143_638 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_142_104 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_108_392 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_43_6 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_150_181 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4020_ _4020_/A1 _4020_/A2 _4020_/A3 _4020_/A4 _4025_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand4_1
XFILLER_29_4 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_37_302 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_64_121 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_37_357 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5971_ _5971_/A1 _7285_/A2 _5987_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_4
XFILLER_92_463 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_64_176 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4922_ input99/Z input98/Z _4922_/A3 _4922_/A4 _4926_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand4_1
X_7710_ _7710_/D _7877_/RN _7726_/CLK _7710_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffsnq_1
XFILLER_92_496 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7641_ _7641_/D _7901_/RN _7864_/CLK _7641_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_60_371 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4853_ _4853_/A1 _7285_/A2 _4857_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_3804_ hold49/Z hold36/Z _3806_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__and2_1
X_4784_ _7515_/Q _7959_/RN _4795_/S VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_4
X_7572_ _7572_/D _7572_/CLK _7572_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_174_741 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_146_421 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3735_ _4380_/B _3734_/Z _3735_/B _7979_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_6523_ hold835/Z _6536_/A2 _6524_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_134_605 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6454_ _6539_/A1 _6468_/A2 _6454_/B _7854_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_161_413 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5405_ _5701_/A2 _5682_/A3 _5405_/B _5406_/C VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_106_318 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_173_295 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6385_ hold854/Z _6400_/A2 _6386_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_142_660 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_5336_ _5394_/A1 _5344_/A2 _5687_/B _5618_/A3 _5337_/C VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor4_1
X_5267_ _5433_/C _5573_/A1 _5722_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_88_747 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_87_224 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_7006_ _7686_/Q _7189_/B1 _7189_/C1 _7654_/Q _7008_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_85_19 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_4218_ _7782_/Q _6299_/A1 _6248_/A1 _7758_/Q _4262_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_5198_ _5015_/B _5371_/C _5197_/Z _7519_/Q _5415_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai31_1
XFILLER_68_460 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_83_430 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4149_ hold38/Z _3881_/Z _4774_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_83_485 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_71_603 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_83_496 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7908_ _7908_/D _7938_/RN _7940_/CLK _7908_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_4
XFILLER_34_34 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_70_179 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_12_747 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_12_736 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_11_202 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_7839_ _7839_/D _7900_/RN _7862_/CLK _7839_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffsnq_1
XFILLER_133_4 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_11_235 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_50_33 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_180_700 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_20_791 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_165_785 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_125_638 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_119_2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_180_744 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_152_446 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_152_457 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_1_2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_133_682 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_120_321 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_78_235 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_78_224 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_182_65 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_94_717 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_115_70 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_94_739 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_19_357 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_46_121 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_74_463 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_34_305 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_46_176 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_47_699 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_34_327 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1250 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_91_73 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_1283 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1272 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1261 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1294 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_116_605 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_11_780 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_143_413 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xhold718 _7843_/Q hold718/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
Xhold707 hold707/I _7690_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
XFILLER_6_250 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xhold729 _7463_/Q hold729/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
XFILLER_124_660 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_124_671 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6170_ _4476_/I _6174_/A2 _6170_/B hold349/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_115_159 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_5121_ _5087_/B _5680_/B2 _5218_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_151_490 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_130_129 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
Xclkbuf_leaf_3_csclk clkbuf_leaf_9_csclk/I _7892_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_34_2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_111_354 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5052_ _5452_/C _5543_/C _5797_/A2 _5064_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor3_2
XFILLER_111_398 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4003_ _7874_/Q _6486_/A1 _4035_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_93_783 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_53_603 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_179_800 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_65_496 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_111_39 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_80_455 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5954_ _5954_/A1 _6537_/A2 _5970_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_4
XFILLER_178_321 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4905_ _5224_/A3 _5224_/A4 _4905_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__and2_1
X_5885_ _4454_/Z _5885_/A2 _5885_/B _7587_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_52_179 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_178_354 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4836_ _7519_/Q _7518_/Q _7520_/Q _7280_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor3_4
XFILLER_139_708 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7624_ _7624_/D _7961_/RN _7624_/CLK _7624_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_178_398 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_7555_ _7555_/D _7314_/Z _4418_/I1 _7555_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffnrnq_1
X_4767_ hold822/Z _4768_/A2 _4768_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_6506_ hold876/Z _6519_/A2 _6507_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_4698_ _4718_/A1 _4698_/A2 _4698_/B _7438_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_107_638 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_106_104 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7486_ _7486_/D _7503_/CLK _7486_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_3718_ _7907_/Q _6634_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__inv_2
XFILLER_174_593 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_162_744 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_106_148 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_3649_ _7903_/Q _6565_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_6437_ _6539_/A1 _6451_/A2 _6437_/B _7846_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_121_107 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_20_69 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6368_ hold665/Z _6383_/A2 _6369_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_5319_ _5563_/B2 _5365_/B1 _5319_/B _5319_/C _5419_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi211_4
XFILLER_102_321 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_437 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
Xhold12 hold12/I hold12/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
X_6299_ _6299_/A1 _6537_/A2 _6315_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_4
Xhold23 hold23/I hold23/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
XFILLER_29_34 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_48_408 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
Xhold45 hold45/I hold45/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
Xhold34 hold34/I hold34/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
Xhold56 hold56/I hold56/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
Xhold67 hold67/I hold67/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
XFILLER_91_709 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xhold89 hold89/I hold89/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
Xhold78 hold78/I hold78/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
XFILLER_17_806 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_56_463 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_28_176 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_45_33 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_44_636 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_300 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_45_77 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_333 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_322 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_311 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_71_499 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_355 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_344 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_169_354 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_157_505 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_61_10 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_12_522 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_169_387 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_138_741 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_106_671 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_3_286 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_126_80 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_121_641 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xclkbuf_3_2__f_wb_clk_i clkbuf_0_wb_clk_i/Z _7940_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_120_162 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_75_783 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_62_433 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_47_496 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_34_179 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_5670_ _5799_/A1 _5799_/A2 _5776_/A4 _5799_/A3 _5671_/A4 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand4_1
XFILLER_96_4 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1091 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1080 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_4621_ _7990_/I _4652_/A1 _4624_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_175_357 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_163_508 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_129_763 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_30_385 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_7340_ _7340_/D _7295_/Z _7972_/CLK _7340_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
X_4552_ hold816/Z _4553_/A2 _4553_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_7271_ _7271_/A1 _7271_/A2 _7272_/C VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
Xhold515 hold515/I _4657_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
XFILLER_144_744 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xhold526 hold526/I _6117_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
Xhold504 hold504/I _6206_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
XFILLER_7_570 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4483_ hold319/Z _4487_/A1 _4487_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_6222_ hold370/Z _6225_/A2 _6223_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
Xhold559 hold559/I _7426_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
Xhold537 hold537/I _6100_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
Xhold548 _7562_/Q hold548/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
XFILLER_143_298 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_106_17 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_103_129 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_103_118 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_103_107 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6153_ _4476_/I _6157_/A2 _6153_/B hold224/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
XTAP_820 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_831 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_842 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_853 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_6084_ hold345/Z _6089_/A2 hold346/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_5104_ _5705_/A2 _5783_/A2 _5104_/B _5105_/A4 VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
XTAP_864 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_875 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_886 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_5035_ _5069_/A2 _4930_/Z _4953_/Z _5035_/A4 _5099_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand4_4
XFILLER_73_709 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_897 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_38_463 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_38_485 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_53_422 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_80_252 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_25_135 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6986_ _6986_/A1 _6986_/A2 _6991_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_179_641 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5937_ _5937_/A1 _7285_/A2 _5953_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_4
XFILLER_40_105 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_53_499 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_40_127 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_7607_ _7607_/D _7961_/RN _7624_/CLK _7607_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffsnq_2
X_5868_ _4454_/Z _5868_/A2 _5868_/B _7580_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_21_352 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5799_ _5799_/A1 _5799_/A2 _5799_/A3 _5799_/A4 _5800_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand4_1
X_4819_ _7219_/A1 _4828_/S _4819_/B _7496_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_31_24 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_135_700 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_5_518 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7538_ _7538_/D _7961_/RN _7650_/CLK _7538_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_147_68 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_147_46 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_134_210 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7469_ _7469_/D _7938_/RN _7639_/CLK _7469_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_150_747 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_212 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
Xinput102 wb_adr_i[16] _4924_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_1
XFILLER_103_641 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xinput124 wb_adr_i[7] _3727_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_12
Xinput113 wb_adr_i[26] _3661_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyb_1
Xinput135 wb_dat_i[16] _7239_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XFILLER_130_471 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_103_696 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_1_779 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
Xinput146 wb_dat_i[26] _7250_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyb_1
Xinput157 wb_dat_i[7] _7277_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XFILLER_102_173 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_56_32 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_63_219 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_29_463 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_72_720 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_29_496 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_29_485 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_44_400 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_56_260 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_56_271 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_57_783 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_71_241 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_16_124 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_44_444 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_112_71 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_16_179 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_31_105 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_44_477 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XPHY_152 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_141 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_130 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_185 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_174 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_163 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_173_806 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_157_357 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_157_368 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_196 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_126_744 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_126_788 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_125_298 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_98_138 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_98_105 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_95_812 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_67_525 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
Xclkbuf_leaf_83_csclk _7407_/CLK _7547_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
X_6840_ _7797_/Q _6893_/A2 _6893_/B1 _7773_/Q _6893_/C1 _7635_/Q _6843_/A1 VDD VSS
+ gf180mcu_fd_sc_mcu7t5v0__aoi222_1
XFILLER_63_753 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
Xclkbuf_leaf_98_csclk _7407_/CLK _7767_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
X_6771_ _6771_/A1 _6771_/A2 _6771_/A3 _6771_/A4 _6777_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand4_1
XFILLER_22_105 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_35_499 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5722_ _5722_/A1 _5620_/B _5722_/B _5723_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_3983_ _7352_/Q hold194/I _4505_/A1 _7368_/Q _3985_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_16_680 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_22_138 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_164_806 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5653_ _5653_/A1 _5542_/Z _5764_/A2 _5746_/A4 _5654_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor4_1
X_5584_ _5704_/A1 _5716_/A2 _5732_/A2 _5794_/A2 _5589_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand4_1
X_4604_ _4604_/A1 _6537_/A2 _4608_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_7323_ _7877_/RN _4334_/Z _7323_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__and2_1
X_4535_ hold895/Z _4548_/A2 _4536_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_144_530 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
Xclkbuf_leaf_36_csclk _7422_/CLK _7852_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
Xhold301 hold301/I _7868_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
XFILLER_7_70 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xhold312 _7635_/Q hold312/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
Xhold323 _7997_/I hold323/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
Xhold334 hold334/I _7689_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
Xhold367 _7596_/Q hold367/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
X_7254_ _7518_/Q _7254_/A2 _7256_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_132_747 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_131_224 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
Xhold378 _7764_/Q hold378/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
Xhold345 _7681_/Q hold345/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
Xhold356 hold356/I _7657_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
X_4466_ _7350_/Q _4487_/A1 _4467_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
Xhold389 _7780_/Q hold389/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
X_4397_ _7438_/Q input58/Z _7335_/Q _4397_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_6205_ hold503/Z _6208_/A2 hold504/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_7185_ _7433_/Q _7938_/Q _7185_/B _7187_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_131_268 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_112_460 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6136_ _4476_/I _6140_/A2 _6136_/B hold337/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_86_812 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_650 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_661 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_672 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_683 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_694 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_58_558 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_6067_ hold326/Z _6072_/A2 hold327/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_5018_ _5529_/A2 _5529_/A3 _5528_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_2
XFILLER_26_24 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_39_783 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1816 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1805 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1849 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1838 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1827 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_26_488 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_53_274 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6969_ _7846_/Q _7193_/A2 _7205_/A2 _7732_/Q _6971_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_167_611 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_10_812 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_158_34 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_158_12 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_155_806 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_139_357 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_21_171 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_21_160 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_42_67 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_182_625 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_166_176 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_158_78 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_127_508 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_108_744 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_108_733 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_5_337 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_101_2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_5_348 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_5_359 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xhold890 _7661_/Q hold890/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
XFILLER_103_460 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_77_812 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_67_97 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_37_709 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_123_70 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_83_30 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_17_444 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_45_753 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_44_263 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_17_499 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_157_176 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_145_316 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_8_131 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_40_491 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_172_179 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4320_ _7336_/Q _4300_/C _4322_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_126_585 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_99_425 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_114_747 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_4_392 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4251_ _7644_/Q _6005_/A1 _4883_/A1 _7533_/Q _4253_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_86_108 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_68_812 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4182_ _7693_/Q _6107_/A1 _4858_/A1 _7524_/Q _4183_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_7941_ _7941_/D _7959_/RN _7959_/CLK _7941_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_103_29 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_94_174 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_82_325 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7872_ _7872_/D _7901_/RN _7872_/CLK _7872_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffsnq_1
XFILLER_36_753 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_51_712 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_90_380 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6823_ _7714_/Q _6885_/B1 _6890_/A2 _7642_/Q _6824_/A4 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_23_425 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_149_611 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3966_ _7673_/Q _6056_/A1 _5937_/A1 _7617_/Q _3992_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_6754_ _6754_/A1 _6767_/C _6754_/B1 _6754_/B2 _7433_/Q _6755_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi221_1
XFILLER_50_266 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_148_121 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_137_806 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5705_ _5104_/B _5705_/A2 _5705_/B _5706_/A4 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_10_108 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_6685_ _7604_/Q _7910_/Q _6879_/A1 _6686_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor3_1
XFILLER_176_463 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_164_614 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_5636_ _5636_/A1 _5417_/I _5708_/B _5679_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor3_1
X_3897_ _7755_/Q _6226_/A1 _6401_/A1 _7837_/Q _3901_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_148_176 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_128_37 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_12_37 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_105_703 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5567_ _4998_/B _5412_/B _5567_/A3 _5706_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor3_1
XFILLER_88_19 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_3_808 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xhold131 _7443_/Q hold131/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
X_5498_ _5689_/A2 _5498_/A2 _5498_/B _5543_/C _5653_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi211_1
X_7306_ _7901_/RN _4334_/Z _7306_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_117_596 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4518_ hold473/Z _4521_/A2 hold474/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
Xhold153 hold153/I _5928_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
XFILLER_2_318 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xhold120 hold120/I _7651_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
Xhold142 hold142/I _4727_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
X_7237_ _7516_/Q _7237_/A2 _7280_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_4449_ hold46/Z _4449_/A2 hold50/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
Xhold186 hold186/I _7683_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
Xhold164 _7793_/Q hold164/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
Xhold175 hold175/I _7761_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
XFILLER_78_609 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_5_9 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
Xhold197 hold197/I _6072_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
XFILLER_120_717 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_59_812 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_132_599 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_113_780 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7168_ _7168_/A1 _7168_/A2 _7178_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_6119_ _4476_/I _6123_/A2 _6119_/B hold331/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_7099_ _7737_/Q _7205_/A2 _7205_/B1 _7745_/Q _7100_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_85_141 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_74_804 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_491 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_480 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_19_709 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_100_463 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2325 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2314 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2303 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_27_753 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_37_89 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2369 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2347 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2358 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2336 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_160_79 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1624 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1613 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1602 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1657 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1646 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1635 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_26_296 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_41_200 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_41_211 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_42_756 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_53_33 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_149_2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1679 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1668 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_53_77 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_53_88 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_6_602 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_182_422 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_139_176 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_10_686 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_154_146 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_6_646 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_154_179 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_150_330 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xclkbuf_1_0__f__1040_ clkbuf_0__1040_/Z _4826_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_68_108 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_49_388 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_91_144 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_64_358 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_91_155 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_33_712 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_178_717 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_150_90 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3820_ hold26/Z _3925_/A2 hold75/Z _3963_/A4 hold76/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand4_4
XFILLER_60_564 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3751_ _3730_/Z _3751_/A2 _3751_/A3 _3752_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor3_1
XFILLER_158_463 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_119_806 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_145_102 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3682_ _7841_/Q _3682_/ZN VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_6470_ hold787/Z _6485_/A2 _6471_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_145_157 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5421_ _5421_/A1 _5421_/A2 _5421_/A3 _5421_/B1 _5498_/A2 _5422_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai32_1
XFILLER_64_2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
Xoutput214 _4411_/Z mgmt_gpio_out[14] VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_1
XFILLER_173_499 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_160_105 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_145_168 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
Xoutput225 _7998_/Z mgmt_gpio_out[24] VDD VSS gf180mcu_fd_sc_mcu7t5v0__buf_4
X_5352_ _5788_/A2 _5534_/A2 _5353_/A4 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_99_211 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
Xoutput203 _3708_/ZN mgmt_gpio_oeb[4] VDD VSS gf180mcu_fd_sc_mcu7t5v0__buf_4
X_4303_ _7414_/Q _4297_/Z _4303_/A3 _4303_/B _4304_/I0 VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai31_1
Xoutput236 _8006_/Z mgmt_gpio_out[34] VDD VSS gf180mcu_fd_sc_mcu7t5v0__buf_4
XFILLER_126_382 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_114_544 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_5_690 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xoutput258 _7567_/Q pll90_sel[1] VDD VSS gf180mcu_fd_sc_mcu7t5v0__buf_4
Xoutput247 _4418_/Z pad_flash_clk VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_1
X_7022_ _7734_/Q _7205_/A2 _7205_/B1 _7742_/Q _7023_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_5283_ _5247_/B _5624_/B _5783_/B _5288_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_87_428 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xoutput269 _7564_/Q pll_sel[1] VDD VSS gf180mcu_fd_sc_mcu7t5v0__buf_4
XFILLER_99_288 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4234_ _7604_/Q _5920_/A1 _4873_/A1 _7529_/Q _4236_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_114_17 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_67_141 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4165_ _7815_/Q _6367_/A1 _4609_/A1 _7408_/Q _4843_/A1 _7508_/Q _4167_/A3 VDD VSS
+ gf180mcu_fd_sc_mcu7t5v0__aoi222_1
XFILLER_56_804 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_4096_ _7377_/Q hold55/I _4239_/A2 input22/Z _4719_/A1 input63/Z _4100_/A1 VDD VSS
+ gf180mcu_fd_sc_mcu7t5v0__aoi222_1
XFILLER_83_667 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7924_ _7924_/D _7938_/RN _4411_/I1 _7924_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_55_369 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_169_706 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_7855_ _7855_/D _7900_/RN _7878_/CLK _7855_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffsnq_1
XFILLER_24_723 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_51_531 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6806_ _7706_/Q _6889_/A2 _6805_/Z _6830_/B _6819_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_4998_ _5705_/A2 _4996_/Z _4998_/B _4998_/C _4999_/A4 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi211_1
X_7786_ _7786_/D _7900_/RN _7892_/CLK _7786_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_11_428 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_177_783 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6737_ _7793_/Q _6893_/A2 _6893_/B1 _7769_/Q _6738_/A4 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_3949_ input59/Z _5886_/A1 _4219_/A2 input18/Z _6469_/A1 _7868_/Q _3953_/A1 VDD VSS
+ gf180mcu_fd_sc_mcu7t5v0__aoi222_2
XFILLER_149_496 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6668_ _7375_/Q _6882_/A2 _6665_/Z _7740_/Q _6683_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_5619_ _5319_/C _5714_/B1 _5319_/B _5619_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__or3_1
X_6599_ _7912_/Q _6599_/A2 _6599_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__or2_4
XFILLER_151_116 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_136_179 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_155_46 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_117_382 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_105_566 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_105_555 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_59_653 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_101_783 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_2100 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_104_72 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_73_144 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_2144 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2133 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2111 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2122 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_15_712 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_34_509 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_2177 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2166 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2155 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1432 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1421 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1410 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_531 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2199 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2188 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1454 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1465 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1443 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1498 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1487 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1476 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_80_64 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_10_450 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_116_809 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_182_274 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_170_403 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_155_499 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_142_138 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_89_73 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_151_661 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_96_203 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_69_406 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_150_160 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_69_428 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_96_247 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_49_141 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_65_667 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_65_645 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5970_ _6553_/A1 _5970_/A2 _5970_/B hold140/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_52_317 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4921_ _4917_/Z _4919_/Z _5210_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_4
XFILLER_64_188 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_33_531 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_100_19 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7640_ _7640_/D _7901_/RN _7858_/CLK _7640_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
X_4852_ _4454_/Z _4852_/A2 _4852_/B _7510_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_3803_ _7341_/Q hold147/Z _7414_/Q _3803_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_7571_ _7571_/D _7961_/RN _7650_/CLK _7571_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffsnq_1
XFILLER_20_247 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_21_759 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_4783_ _4454_/Z _4783_/A2 _4783_/B _7477_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_159_783 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3734_ _7414_/Q _7413_/Q _7411_/Q _3734_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__or3_2
XFILLER_146_400 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_118_102 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_20_269 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6522_ _6539_/A1 _6536_/A2 _6522_/B _7886_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_3665_ _7607_/Q _6754_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_6453_ hold799/Z _6468_/A2 _6454_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_9_292 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_161_425 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5404_ _5404_/A1 _5779_/B1 _5682_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_133_116 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_118_179 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_133_138 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6384_ _6384_/A1 hold5/Z _6400_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_4
XFILLER_142_672 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_142_650 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_130_812 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5335_ _5335_/A1 _5335_/A2 _5331_/Z _5335_/A4 _5354_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand4_1
XFILLER_126_190 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5266_ _5687_/B _5645_/A3 _5680_/B1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_114_385 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_114_396 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7005_ _7678_/Q _7191_/A2 _7190_/B1 _7614_/Q _7190_/A2 _7792_/Q _7008_/A2 VDD VSS
+ gf180mcu_fd_sc_mcu7t5v0__aoi222_1
X_4217_ hold609/Z _4217_/A2 _5871_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_5197_ _5209_/A2 _5209_/A3 _5197_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_56_612 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_110_580 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4148_ hold38/Z _3963_/Z _4764_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_4079_ _7662_/Q _6039_/A1 _6452_/A1 _7856_/Q _4080_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_18_69 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_55_144 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_70_114 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7907_ _7907_/D _7938_/RN _7938_/CLK _7907_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffsnq_4
XFILLER_24_531 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_51_361 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7838_ _7838_/D _7900_/RN _7862_/CLK _7838_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffsnq_1
XFILLER_157_709 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7769_ _7769_/D _7900_/RN _7897_/CLK _7769_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_109_113 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_166_34 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_109_124 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_137_499 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_121_812 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_59_32 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_105_396 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xclkbuf_3_1__f_wb_clk_i clkbuf_0_wb_clk_i/Z _7949_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_78_247 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_59_87 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_182_99 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_120_388 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_94_729 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_101_591 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_101_580 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_46_188 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_131_70 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_131_81 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1240 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_91_52 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1284 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1273 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1262 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1251 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_372 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1295 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_30_534 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_156_731 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_171_712 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xhold719 _7851_/Q hold719/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
Xhold708 _7618_/Q hold708/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
XFILLER_7_763 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_115_138 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_6_273 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_130_108 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_124_650 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_112_812 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5120_ _5319_/C _5689_/A2 _5390_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_5051_ _5006_/C _5448_/A1 _5797_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_4
XFILLER_97_567 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_85_707 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_27_2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4002_ _4002_/A1 _4427_/B _4002_/B1 _4002_/B2 _7553_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_37_100 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_38_656 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_92_250 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_65_453 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_1_83 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_25_306 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_37_144 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_37_188 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_179_812 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5953_ _6553_/A1 _5953_/A2 _5953_/B hold138/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_4904_ _5087_/C _4900_/Z _5496_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_4
X_5884_ hold862/Z _5885_/A2 _5885_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_52_169 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4835_ _4454_/Z _4835_/A2 _4835_/B _7505_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_7623_ hold77/Z _7961_/RN _7960_/CLK _7623_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_147_731 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_4766_ _6539_/A1 _4768_/A2 _4766_/B _7470_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_21_567 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7554_ _7554_/D _7313_/Z _4418_/I1 _7554_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffnrnq_1
X_6505_ _6539_/A1 _6519_/A2 _6505_/B _7878_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_3717_ _7910_/Q _6878_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_12
XFILLER_146_263 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4697_ hold491/Z _3819_/Z _4697_/B _4698_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_119_477 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_119_488 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7485_ _7485_/D _7949_/CLK _7485_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_162_756 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_119_499 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6436_ hold795/Z _6451_/A2 _6437_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_20_37 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_3648_ _7432_/Q _6572_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_136_59 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_136_48 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_136_37 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_122_609 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6367_ _6367_/A1 _7285_/A2 _6383_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_4
X_5318_ _5350_/A3 _5495_/B2 _5555_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_2
XFILLER_88_534 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xhold13 hold13/I hold13/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
XFILLER_130_653 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6298_ _6553_/A1 _6298_/A2 _6298_/B _7781_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_88_567 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xhold35 hold35/I hold35/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
Xhold46 hold46/I hold46/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
X_5249_ _3728_/I _5022_/B _5054_/Z _5687_/B _5425_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor4_4
Xhold24 hold24/I hold24/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
Xhold57 hold57/I hold57/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
Xhold68 hold68/I hold68/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
Xhold79 hold79/I hold79/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
XFILLER_68_291 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_56_442 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_84_795 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_83_283 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_301 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_169_311 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_334 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_323 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_312 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_356 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_345 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_169_366 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_157_517 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_101_84 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_101_73 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_12_534 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_24_383 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_131_2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_8_516 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_138_731 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_165_550 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_153_712 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_6_17 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_180_531 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_152_211 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_152_200 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_125_436 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_125_425 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_4_744 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_121_620 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_112_108 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_105_160 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_79_512 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_121_631 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_79_567 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_66_239 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_74_250 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_19_144 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_142_91 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_35_659 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1092 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1081 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1070 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_30_331 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4620_ _4620_/A1 _5903_/A2 _4686_/B1 _3830_/Z hold22/Z _4652_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi221_4
XFILLER_129_720 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4551_ _6539_/A1 _4553_/A2 _4551_/B _7383_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_7270_ _7520_/Q _7270_/A2 _7270_/B1 _7518_/Q _7271_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_1
Xhold516 hold516/I _7424_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
XFILLER_144_756 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xhold527 hold527/I _7696_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
Xhold505 hold505/I _7738_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
X_4482_ _4487_/A1 _4481_/I _4482_/B _7353_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_6221_ _4476_/I _6225_/A2 _6221_/B hold339/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
Xhold538 hold538/I _7688_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
XFILLER_104_609 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_89_309 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
Xhold549 _7614_/Q hold549/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
X_6152_ hold222/Z _6157_/A2 hold223/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_131_428 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_810 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_106_29 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5103_ _5669_/B _5669_/A1 _5648_/A2 _5104_/B _5105_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XTAP_821 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_832 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_843 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_111_141 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_100_804 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_6083_ _6547_/A1 _6089_/A2 _6083_/B hold544/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
XTAP_854 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_865 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_876 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_5034_ _5661_/A1 _4965_/B _5647_/A2 _5752_/B1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor3_4
XFILLER_66_740 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_887 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_898 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_122_17 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_93_570 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_93_581 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_65_283 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6985_ _7693_/Q _7194_/A2 _7194_/B1 _7661_/Q _7194_/C1 _7807_/Q _6986_/A2 VDD VSS
+ gf180mcu_fd_sc_mcu7t5v0__aoi222_1
X_5936_ _6553_/A1 _5936_/A2 _5936_/B hold206/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_40_117 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_178_163 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_166_325 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5867_ hold765/Z _5868_/A2 _5868_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_7606_ _7606_/D _7961_/RN _7606_/CLK _7606_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_182_807 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5798_ _5583_/C _5185_/B _5798_/A3 _5798_/A4 _5799_/A4 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor4_1
X_4818_ _7496_/Q _4828_/S _4819_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_4749_ hold418/Z _4749_/I1 _4753_/S _4749_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_135_712 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7537_ _7537_/D _7961_/RN _7650_/CLK _7537_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_162_531 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_107_425 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7468_ _7468_/D _7961_/RN _7639_/CLK _7468_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_134_266 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6419_ hold789/Z _6434_/A2 _6420_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_122_417 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_89_810 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7399_ _7399_/D input75/Z _7477_/CLK _7399_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
Xinput114 wb_adr_i[27] _4368_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyb_1
Xinput125 wb_adr_i[8] _4923_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyb_1
Xinput103 wb_adr_i[17] _4924_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyb_1
Xinput136 wb_dat_i[17] _7244_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XFILLER_76_504 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_279 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xinput158 wb_dat_i[8] _7240_/B1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyb_1
Xinput147 wb_dat_i[27] _7255_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XFILLER_102_196 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_76_548 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_179_2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_29_475 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_56_250 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_72_743 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_72_32 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_13_810 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_44_467 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_169_141 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_71_286 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_142 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_131 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_120 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_157_314 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_175 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_164 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_153 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
Xclkbuf_leaf_2_csclk clkbuf_leaf_9_csclk/I _7887_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XPHY_197 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_186 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_12_375 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_8_313 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_40_673 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_145_509 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_113_428 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_98_128 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_180_394 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_140_258 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_140_247 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_97_73 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_39_239 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_94_389 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_75_570 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_47_283 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3982_ _7851_/Q _6435_/A1 _6469_/A1 _7867_/Q _3985_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_6770_ _7818_/Q _6880_/A2 _6893_/C1 _7632_/Q _6771_/A4 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_63_798 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XPHY_0 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
X_5721_ _5621_/B _5724_/A2 _5721_/B _5721_/C _5722_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XFILLER_94_2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_176_601 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_31_651 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_50_459 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5652_ _5162_/B _5652_/A2 _5652_/A3 _5652_/A4 _5746_/A4 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand4_1
XFILLER_30_172 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_175_177 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_175_144 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_117_712 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5583_ _5062_/Z _5690_/A1 _5583_/B _5583_/C _5794_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi211_1
X_4603_ _4454_/Z _4603_/A2 _4603_/B _7404_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_7322_ _7877_/RN _4334_/Z _7322_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__and2_1
X_4534_ _6539_/A1 _4548_/A2 _4534_/B _7375_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
Xhold302 _7715_/Q hold302/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
XFILLER_116_211 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
Xhold324 hold324/I _4652_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
XFILLER_144_542 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
Xhold313 _7813_/Q hold313/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
Xhold335 _7705_/Q hold335/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
XFILLER_7_93 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_7253_ _7253_/A1 _7277_/B _7253_/B _7952_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi21_1
Xhold368 hold368/I _5905_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
X_4465_ hold64/I _4748_/I1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
Xhold346 hold346/I _6085_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
XFILLER_116_277 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xhold357 _7370_/Q hold357/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
Xhold379 hold379/I _6262_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
X_6204_ _4476_/I _6208_/A2 _6204_/B hold352/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_4396_ _7447_/Q input81/Z _4396_/S _4396_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_7184_ _7184_/A1 _7210_/A2 _7184_/B1 _7184_/B2 _7433_/Q _7185_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi221_1
X_6135_ hold335/Z _6140_/A2 hold336/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_98_673 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_640 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_651 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_6066_ _6547_/A1 _6072_/A2 _6066_/B hold547/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_85_323 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_662 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_673 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_684 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_695 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_58_548 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5017_ _5230_/A1 _5024_/A2 _5200_/B _5529_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_4
XFILLER_38_250 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_39_773 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1806 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1839 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1828 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1817 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_26_478 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_26_467 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6968_ _7758_/Q _7202_/C2 _7201_/A2 _7748_/Q _6971_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_53_286 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5919_ hold2/Z _5919_/A2 hold9/Z hold10/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_10_802 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_6899_ _7930_/Q _7133_/S _6900_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_22_662 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_6_806 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_107_200 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_107_211 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_181_169 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_108_756 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_174_45 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_174_34 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_162_383 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_150_534 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_122_247 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xhold891 _7526_/Q hold891/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
Xhold880 _7847_/Q hold880/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
XFILLER_107_61 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_89_651 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_88_194 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_76_356 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_123_60 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_76_389 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_57_570 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_123_93 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_72_540 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_29_283 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_17_489 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_45_798 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_72_584 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_158_601 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_9_611 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_32_459 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_173_615 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_157_144 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_145_306 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_173_637 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_172_125 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_9_699 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_8_176 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_126_531 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_153_361 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_113_225 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_4250_ _7620_/Q _5954_/A1 _4812_/A1 _7494_/Q _4253_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_141_567 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_68_802 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4181_ _7733_/Q _6192_/A1 _4878_/A1 _7532_/Q _4868_/A1 _7528_/Q _4183_/A2 VDD VSS
+ gf180mcu_fd_sc_mcu7t5v0__aoi222_1
X_7940_ _7940_/D _7961_/RN _7940_/CLK _7940_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
X_7871_ _7871_/D _7875_/RN _7874_/CLK _7871_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffsnq_1
X_6822_ _7722_/Q _6881_/A2 _6881_/B1 _7698_/Q _6824_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_36_798 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_90_392 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_35_286 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6753_ _6753_/A1 _6753_/A2 _6753_/A3 _6754_/B2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor3_1
XFILLER_51_779 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3965_ _7649_/Q _6005_/A1 _4231_/B1 input68/Z _3994_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_176_420 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_149_634 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_148_133 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_148_100 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3896_ _3896_/A1 _3896_/A2 _3896_/A3 _3918_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand3_2
X_5704_ _5704_/A1 _5704_/A2 _5704_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__and2_1
X_6684_ _6684_/A1 _6684_/A2 _6684_/A3 _6686_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor3_1
XFILLER_148_166 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5635_ _5692_/B _5218_/C _5708_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_1
Xhold110 _7687_/Q hold110/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
XFILLER_117_542 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5566_ _5602_/A2 _4993_/B _5663_/A1 _5566_/B _5567_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai31_1
Xhold132 hold132/I _4718_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
XFILLER_172_670 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5497_ _5452_/C _5498_/A2 _5497_/A3 _5499_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor3_1
X_7305_ _7901_/RN _4334_/Z _7305_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__and2_1
Xhold121 _7695_/Q hold121/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
X_4517_ _6549_/A1 _4521_/A2 _4517_/B hold744/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
Xhold143 hold143/I _7447_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
X_7236_ _3658_/I _7236_/A2 _7237_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_4448_ hold46/Z _4449_/A2 hold47/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__and2_4
XFILLER_132_534 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xhold165 hold165/I _6324_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
XFILLER_104_247 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xhold176 _7897_/Q hold176/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
Xhold154 hold154/I _7607_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
XFILLER_144_37 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_144_48 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
Xhold198 hold198/I _7675_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
Xhold187 _7691_/Q hold187/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
XFILLER_59_802 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4379_ _4379_/I _7412_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_7167_ _7509_/Q _7191_/A2 _7190_/B1 _7468_/Q _7190_/A2 _7401_/Q _7168_/A2 VDD VSS
+ gf180mcu_fd_sc_mcu7t5v0__aoi222_1
X_6118_ hold329/Z _6123_/A2 hold330/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_7098_ _7779_/Q _7200_/A2 _7200_/B1 _7867_/Q _7100_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_86_676 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_492 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_481 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_470 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_58_356 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6049_ hold16/Z _6055_/A2 _6049_/B hold39/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_37_35 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_39_570 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_58_389 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2326 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2315 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2304 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_170_6 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2348 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2359 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2337 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1614 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1603 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_702 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1658 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1647 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1636 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1625 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1669 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_41_256 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_179_280 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_182_401 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_139_166 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_139_144 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xclkbuf_leaf_82_csclk clkbuf_leaf_9_csclk/I _7790_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_154_114 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_108_520 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_10_676 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_154_136 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_108_531 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_182_489 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_182_478 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xclkbuf_leaf_97_csclk _7407_/CLK _7881_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_135_383 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_123_545 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_7917__361 _7917_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__tieh
XFILLER_123_567 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_111_718 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xclkbuf_leaf_20_csclk _7873_/CLK _7896_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_92_635 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_92_602 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_49_378 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_91_134 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_18_721 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
Xclkbuf_leaf_35_csclk _7422_/CLK _7812_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_17_231 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_150_80 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_72_392 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_17_286 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_60_554 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3750_ _7411_/Q _3774_/A2 _3751_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_20_429 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_32_267 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_173_423 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3681_ _7849_/Q _3681_/ZN VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_5420_ _5062_/Z _5176_/B _5421_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_9_496 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xoutput215 _4410_/Z mgmt_gpio_out[15] VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_1
X_5351_ _5498_/A2 _5622_/A1 _5534_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_1
Xoutput226 _7999_/Z mgmt_gpio_out[25] VDD VSS gf180mcu_fd_sc_mcu7t5v0__buf_4
XFILLER_99_201 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xoutput204 _3707_/ZN mgmt_gpio_oeb[5] VDD VSS gf180mcu_fd_sc_mcu7t5v0__buf_4
XFILLER_57_2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
Xoutput237 _4396_/Z mgmt_gpio_out[35] VDD VSS gf180mcu_fd_sc_mcu7t5v0__buf_4
X_4302_ _4308_/S _4296_/Z _7342_/Q _4303_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_114_534 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5282_ _5282_/A1 _5282_/A2 _5282_/A3 _5298_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand3_1
Xoutput259 _7568_/Q pll90_sel[2] VDD VSS gf180mcu_fd_sc_mcu7t5v0__buf_4
Xoutput248 _4436_/Z pad_flash_clk_oe VDD VSS gf180mcu_fd_sc_mcu7t5v0__buf_4
XFILLER_141_353 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_102_729 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7021_ _7824_/Q _7202_/A2 _7204_/B1 _7768_/Q _7025_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_4233_ _7375_/Q hold55/I hold43/I _7740_/Q _4256_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_4164_ _7400_/Q _4589_/A1 _4527_/A1 _7374_/Q _4167_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_4095_ _7888_/Q _6520_/A1 hold43/I _7742_/Q _4106_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_68_676 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_67_164 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_7923_ _7923_/D _7923_/RN _4411_/I1 _7923_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_55_359 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_70_318 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_130_28 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7854_ _7854_/D _7901_/RN _7854_/CLK _7854_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffsnq_1
XFILLER_23_212 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_168_206 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_7785_ _7785_/D _7900_/RN _7897_/CLK _7785_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
X_6805_ _7738_/Q _6878_/A2 _6805_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__or2_1
X_4997_ _3722_/I _3723_/I _5006_/B _5006_/C _5663_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand4_4
XFILLER_149_420 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6736_ _7825_/Q _6891_/A2 _6891_/B1 _7671_/Q _6891_/C1 _7777_/Q _6738_/A3 VDD VSS
+ gf180mcu_fd_sc_mcu7t5v0__aoi222_1
XFILLER_176_250 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_149_442 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_3948_ _3948_/A1 _3948_/A2 _3948_/A3 _3948_/A4 _3954_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand4_2
XFILLER_176_261 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_137_637 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_136_103 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3879_ hold609/Z _3869_/I _3879_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__or2_4
XFILLER_109_339 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_99_19 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_6667_ _7684_/Q _6884_/B1 _6892_/B1 _7724_/Q _6681_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_5618_ _5689_/A1 _5692_/B _5618_/A3 _5618_/B1 _5620_/B _5632_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai32_1
X_6598_ _7434_/Q _7912_/Q _7911_/Q _6609_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_133_810 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5549_ _5765_/A2 _5803_/A4 _5549_/A3 _5765_/A3 _5557_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand4_1
XFILLER_117_361 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_105_512 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_155_58 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_2_105 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xclkbuf_3_0__f_wb_clk_i clkbuf_0_wb_clk_i/Z _7503_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_160_673 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_160_695 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_7219_ _7219_/A1 _7228_/S _7219_/B _7942_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_48_34 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_171_35 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_100_250 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_86_484 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_74_602 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_74_613 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2101 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_104_51 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_104_62 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_86_495 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_19 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_58_197 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2134 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2112 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2123 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_73_156 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_27_540 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_27_551 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_27_562 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2167 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2156 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_161_2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2145 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1433 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1422 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1411 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1400 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2189 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2178 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_120_50 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1455 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1466 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1444 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_9_17 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_54_392 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_159_239 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1499 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1488 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1477 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_14_267 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_80_43 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_167_283 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_128_648 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_13_70 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_129_70 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_124_810 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_89_30 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_182_297 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_170_459 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_89_85 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_150_194 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_145_91 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_96_259 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_49_131 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_65_602 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_77_495 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_64_112 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_80_605 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4920_ _4917_/Z _4919_/Z _4920_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__and2_4
XFILLER_178_504 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4851_ hold818/Z _4852_/A2 _4852_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_3802_ _7341_/Q _4383_/A1 _4306_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_4782_ hold834/Z _4783_/A2 _4783_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_21_749 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7570_ _7570_/D _7961_/RN _7570_/CLK _7570_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffsnq_1
XFILLER_158_250 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_158_261 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_146_423 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3733_ _4424_/A1 _3731_/Z _3733_/B _7980_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_119_637 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_20_259 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6521_ hold785/Z _6536_/A2 _6522_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_6452_ _6452_/A1 _6537_/A2 _6468_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_4
X_3664_ _3664_/I _4425_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_5403_ _5579_/B _5591_/A2 _5559_/A1 _5577_/C _5407_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor4_1
XFILLER_118_158 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_115_810 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_173_286 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6383_ _6553_/A1 _6383_/A2 _6383_/B hold159/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_133_128 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5334_ _5404_/A1 _5424_/A1 _5292_/B _5087_/B _5334_/C _5335_/A4 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi221_1
XFILLER_141_161 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_141_150 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_88_738 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_87_215 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5265_ _5624_/A1 _5759_/A1 _5724_/B _5561_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_5196_ _5011_/B _3723_/I _5211_/A3 _4920_/Z _5209_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand4_2
X_7004_ _7702_/Q _7190_/C1 _7008_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_4216_ hold27/I _4075_/B _4238_/B1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_4147_ hold38/Z _4151_/A2 _4779_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_56_602 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_18_37 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_4078_ _7670_/Q _6056_/A1 _5920_/A1 _7606_/Q _4219_/A2 input13/Z _4080_/A2 VDD VSS
+ gf180mcu_fd_sc_mcu7t5v0__aoi222_1
XFILLER_71_638 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7906_ _7906_/D _7938_/RN _7938_/CLK _7906_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_2
X_7837_ _7837_/D _7901_/RN _7869_/CLK _7837_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_36_392 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_169_559 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_34_58 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_7768_ _7768_/D _7901_/RN _7864_/CLK _7768_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffsnq_1
XFILLER_11_215 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_177_570 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7699_ _7699_/D _7923_/RN _7720_/CLK _7699_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
X_6719_ _7614_/Q _6647_/Z _6890_/A2 _7638_/Q _6720_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_149_283 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_50_46 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_137_489 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_109_169 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_152_448 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_3_425 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_121_802 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_105_353 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_79_716 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_3_469 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_1_4 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_182_34 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_78_226 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_47_602 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_101_570 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_87_793 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_75_32 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_62_605 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_35_808 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_131_60 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_34_318 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1241 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1230 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1274 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1263 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1252 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1296 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1285 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_168_581 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_156_798 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_128_467 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
Xhold709 _7875_/Q hold709/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
XFILLER_155_286 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_171_779 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_124_673 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_123_161 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_111_312 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_97_513 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_69_215 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_5050_ _5006_/C _5448_/A1 _5179_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__and2_4
XFILLER_38_602 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4001_ hold949/Z _4284_/A1 _4427_/B _4002_/B2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_77_292 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_93_763 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_1_73 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5952_ hold137/Z _5953_/A2 _5953_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_111_19 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_53_638 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4903_ _3723_/I _4946_/A1 _5648_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_4
XFILLER_18_392 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_52_159 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_178_334 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_80_479 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_61_660 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5883_ _6539_/A1 _5885_/A2 _5883_/B _7586_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_4834_ hold837/Z _4835_/A2 _4835_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_7622_ _7622_/D _7961_/RN _7960_/CLK _7622_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffsnq_1
XFILLER_178_389 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_166_518 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_159_570 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_147_721 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4765_ hold739/Z _4768_/A2 _4766_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_21_557 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7553_ _7553_/D _7312_/Z _4418_/I1 _7553_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffnrnq_1
X_6504_ hold805/Z _6519_/A2 _6505_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_3716_ _7467_/Q _7210_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_4696_ _3819_/Z _4460_/Z _4697_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_7484_ _7484_/D _7949_/CLK _7484_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_3647_ _7511_/Q _7214_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_161_212 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6435_ _6435_/A1 hold5/Z _6451_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_4
XFILLER_161_234 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6366_ _6553_/A1 _6366_/A2 _6366_/B _7813_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_103_802 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5317_ _5768_/A2 _5237_/Z _5624_/B _5648_/B2 _5326_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_1
Xhold14 hold14/I hold14/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
X_6297_ hold258/Z _6298_/A2 _6298_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_152_37 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_152_26 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
Xhold25 hold25/I hold25/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
XFILLER_130_676 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5248_ _5338_/A1 _5369_/B _5303_/A3 _5618_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand3_4
Xhold36 hold36/I hold36/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
Xhold47 hold47/I hold47/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
Xhold58 hold58/I hold58/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
Xhold69 hold69/I hold69/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
X_5179_ _5608_/B _5752_/B1 _5793_/A2 _5179_/B _5188_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai31_1
XFILLER_102_389 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_28_134 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_44_605 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_16_318 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_16_329 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_45_35 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_44_638 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_45_79 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_324 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_313 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_302 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_101_30 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_357 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_346 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_335 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_51_170 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_52_682 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_124_2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_137_286 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_4_756 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_106_673 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_126_60 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_67_708 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_126_93 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_59_270 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_90_733 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_62_413 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_35_638 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_90_744 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_90_799 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_90_788 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_70_490 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1082 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1071 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1060 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_15_373 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_30_321 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1093 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_7_550 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4550_ hold741/Z _4553_/A2 _4551_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
Xhold506 _7441_/Q hold506/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
X_4481_ _4481_/I _4740_/I1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_143_212 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_129_798 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
Xhold517 _7359_/Q hold517/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
X_6220_ hold338/Z _6225_/A2 _6221_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
Xhold528 _7818_/Q hold528/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
XFILLER_116_459 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
Xhold539 _7608_/Q hold539/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
XFILLER_171_576 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6151_ _6547_/A1 _6157_/A2 _6151_/B hold602/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_131_407 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_800 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_5102_ _5669_/A1 _5648_/A2 _5102_/B1 _5777_/A2 _5105_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_106_19 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_811 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_822 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_833 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_844 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_112_676 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_97_354 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6082_ hold542/Z _6089_/A2 hold543/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_855 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_866 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_877 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_5033_ _5199_/B _5201_/B _5369_/B _4944_/Z _5035_/A4 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor4_4
XFILLER_66_730 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_888 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_899 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_26_605 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_81_722 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_6984_ _7847_/Q _7193_/A2 _7193_/B1 _7629_/Q _7193_/C1 _7725_/Q _6986_/A1 VDD VSS
+ gf180mcu_fd_sc_mcu7t5v0__aoi222_1
XFILLER_25_148 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5935_ hold204/Z _5936_/A2 hold205/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_81_799 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_22_800 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_34_671 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5866_ _4481_/I _5868_/A2 _5866_/B _7579_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_21_310 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4817_ _7514_/Q _7959_/RN _4828_/S VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_4
XFILLER_21_354 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7605_ _7605_/D _7961_/RN _7639_/CLK _7605_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
X_5797_ _5797_/A1 _5797_/A2 _5797_/B _5797_/C _5798_/A4 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XFILLER_181_318 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4748_ hold464/Z _4748_/I1 _4753_/S _7461_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_7536_ _7536_/D _7900_/RN _7823_/CLK _7536_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_174_381 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_174_392 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4679_ _3879_/Z _4481_/I _4680_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_134_212 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_119_286 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_7467_ _7467_/D _7900_/RN _7767_/CLK _7467_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_162_543 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_135_779 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6418_ _6418_/A1 hold5/Z _6434_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_4
X_7398_ _7398_/D _7875_/RN _7823_/CLK _7398_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
X_6349_ _6553_/A1 _6349_/A2 _6349_/B hold203/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_88_321 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
Xinput126 wb_adr_i[9] _4925_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyc_1
Xinput115 wb_adr_i[28] _4368_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XFILLER_163_69 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
Xinput104 wb_adr_i[18] _4924_/A4 VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_1
XFILLER_0_247 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
Xinput148 wb_dat_i[28] _7260_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyb_1
Xinput159 wb_dat_i[9] _7245_/B1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyb_1
Xinput137 wb_dat_i[18] _7250_/B1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XFILLER_102_164 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_88_387 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_29_421 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_56_34 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_84_560 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_17_638 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_56_262 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_71_232 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_143 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_132 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_121 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_12_321 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_110 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_157_304 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_176 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_165 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_154 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_8_303 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_157_359 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_198 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_187 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_12_387 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_172_318 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_8_347 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_125_212 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_4_531 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_21_70 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_141_716 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_141_727 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_137_70 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_4_575 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_97_85 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_79_354 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3981_ _3981_/A1 _3981_/A2 _3981_/A3 _3990_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_63_777 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_62_254 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_23_619 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5720_ hold80/I _5520_/C _5738_/C VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_31_641 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_176_657 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_176_646 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5651_ _5651_/A1 _5503_/C _5651_/A3 _5651_/A4 _5651_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__and4_1
XFILLER_87_2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5582_ _5578_/Z _5710_/A1 _5582_/A3 _5582_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__and3_1
XFILLER_117_702 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4602_ hold858/Z _4603_/A2 _4603_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_7321_ _7877_/RN _4334_/Z _7321_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_163_318 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4533_ hold864/Z _4548_/A2 _4534_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_7252_ _7252_/A1 _7280_/A2 _7277_/B _7252_/C _7253_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XFILLER_156_392 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xhold325 hold325/I _7423_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
Xhold303 hold303/I _6157_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
Xhold314 _7853_/Q hold314/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
XFILLER_117_779 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4464_ hold62/Z hold49/Z _4464_/B hold63/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_4
Xhold369 hold369/I _7596_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
XFILLER_144_598 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_131_215 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xhold347 hold347/I _7681_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
Xhold336 hold336/I _6136_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
X_6203_ hold350/Z _6208_/A2 hold351/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
Xhold358 hold358/I _4521_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
XFILLER_171_384 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4395_ _7445_/Q input78/Z _4396_/S _4395_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_7183_ _7210_/A2 _7183_/A2 _7183_/A3 _7184_/B2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor3_1
XFILLER_100_602 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_97_140 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6134_ _6547_/A1 _6140_/A2 _6134_/B hold552/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
XTAP_630 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_641 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_652 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_6065_ hold545/Z _6072_/A2 hold546/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_663 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_674 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_685 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_5016_ _5016_/A1 _5016_/A2 _5016_/B _5452_/C VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_4
XFILLER_85_357 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_696 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1807 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_93_390 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_26_37 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_53_221 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_54_733 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_54_744 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1829 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1818 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_6967_ _6967_/A1 _6967_/A2 _6967_/A3 _6977_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand3_1
X_5918_ hold8/Z _5919_/A2 hold9/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_81_585 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6898_ _7433_/Q _7929_/Q _6898_/B1 _6898_/B2 _6900_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_167_657 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_167_635 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5849_ _7961_/RN _5849_/A2 _7285_/A2 _5851_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_21_140 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_167_668 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7519_ _7519_/D _7959_/RN _7959_/CLK _7519_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_4
XFILLER_154_318 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_101_4 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_89_641 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xhold870 _7559_/Q hold870/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
Xhold881 _7621_/Q hold881/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
XFILLER_3_19 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_122_259 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_107_73 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_88_140 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_1_567 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xhold892 hold892/I _4867_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
XFILLER_76_313 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_60_747 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_32_427 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_13_641 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_158_646 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_157_101 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_40_460 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_157_156 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_12_195 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_138_392 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_141_513 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_99_416 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_113_215 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_99_438 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4180_ _7685_/Q _6090_/A1 _4883_/A1 _7534_/Q _4893_/A1 _7538_/Q _4183_/A1 VDD VSS
+ gf180mcu_fd_sc_mcu7t5v0__aoi222_1
XFILLER_94_132 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_67_357 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_94_176 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_82_316 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_63_530 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_7870_ _7870_/D _7961_/RN _7876_/CLK _7870_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffsnq_1
XFILLER_36_744 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6821_ _7658_/Q _6882_/B1 _6647_/Z _7618_/Q _6824_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_23_405 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_90_382 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6752_ _6752_/A1 _6752_/A2 _6752_/A3 _6752_/A4 _6753_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand4_1
XFILLER_50_235 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_50_246 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3964_ hold149/Z _3963_/Z hold150/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_4
X_5703_ _5104_/B _5658_/B _5685_/B _5247_/B _5703_/C _5704_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi221_1
X_3895_ input33/Z _4249_/A2 _4219_/A2 input19/Z _3896_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_6683_ _6683_/A1 _6683_/A2 _6683_/A3 _6683_/A4 _6684_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand4_1
XFILLER_164_605 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5634_ _5790_/A1 _5726_/A1 _5634_/A3 _5634_/A4 _5637_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor4_1
XFILLER_31_482 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_136_318 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7304_ _7901_/RN _4334_/Z _7304_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__and2_1
X_5565_ _5565_/A1 _5565_/A2 _5565_/A3 _5565_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__or3_1
Xhold100 hold100/I _7865_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
Xhold133 hold133/I _7443_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
Xhold111 hold111/I _6098_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
X_5496_ _5496_/A1 _4993_/B _5647_/A2 _5496_/B _5506_/C VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai31_1
Xhold122 hold122/I _6115_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
X_4516_ hold742/Z _4521_/A2 hold743/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
Xhold144 _7881_/Q hold144/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
X_7235_ _7519_/Q _7235_/A2 _7238_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_4447_ input58/Z _3810_/S _4449_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
Xhold155 _7723_/Q hold155/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
Xhold166 hold166/I _7793_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
Xhold177 hold177/I _6545_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
Xhold188 hold188/I _6106_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
XFILLER_113_760 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
Xhold199 _7699_/Q hold199/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
X_7166_ _7166_/A1 _7166_/A2 _7166_/A3 _7183_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand3_1
X_4378_ _7964_/Q _4378_/A2 _4378_/B _4379_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_6117_ _6547_/A1 _6123_/A2 _6117_/B hold527/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_98_460 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_460 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
Xclkbuf_leaf_1_csclk clkbuf_leaf_9_csclk/I _7900_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
X_7097_ _7097_/A1 _7097_/A2 _7097_/A3 _7097_/A4 _7106_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand4_1
XTAP_493 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_482 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_471 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_6048_ _7664_/Q _6055_/A2 _6049_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_2316 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2305 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_160_37 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2349 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2338 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2327 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1615 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1604 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_27_788 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_27_777 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1648 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1637 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1626 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_7999_ _7999_/I _7999_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_42_747 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_53_35 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_169_35 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1659 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_53_79 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_139_101 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_22_460 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_167_443 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_155_638 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_182_457 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_151_800 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_150_321 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_2_810 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_111_708 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_89_460 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_49_357 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_94_31 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_92_614 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_76_176 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_45_530 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_33_725 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_45_574 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_158_410 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_146_605 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_41_780 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_41_791 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_118_318 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_118_329 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3680_ _7857_/Q _3680_/ZN VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_9_486 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_145_137 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_139_690 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_64_4 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xoutput216 _7990_/Z mgmt_gpio_out[16] VDD VSS gf180mcu_fd_sc_mcu7t5v0__buf_4
XFILLER_145_159 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_126_340 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5350_ _5689_/A2 _5687_/B _5350_/A3 _5788_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor3_1
Xoutput205 _3706_/ZN mgmt_gpio_oeb[6] VDD VSS gf180mcu_fd_sc_mcu7t5v0__buf_4
Xoutput238 _4387_/Z mgmt_gpio_out[36] VDD VSS gf180mcu_fd_sc_mcu7t5v0__buf_4
X_4301_ _4301_/A1 _4301_/A2 _7343_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
Xoutput227 _8000_/Z mgmt_gpio_out[26] VDD VSS gf180mcu_fd_sc_mcu7t5v0__buf_4
XFILLER_99_224 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5281_ _5685_/B _5292_/B _5585_/C _5282_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi21_1
Xoutput249 _4417_/Z pad_flash_csb VDD VSS gf180mcu_fd_sc_mcu7t5v0__buf_4
X_7020_ _7760_/Q _7202_/C2 _7202_/B1 _7784_/Q _7025_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_4232_ input34/Z _4232_/A2 _4848_/A1 _7509_/Q _4260_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_141_387 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_99_279 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4163_ _7376_/Q hold55/I _6452_/A1 _7855_/Q _7584_/Q _5874_/A1 _4167_/A1 VDD VSS
+ gf180mcu_fd_sc_mcu7t5v0__aoi222_1
X_4094_ _7760_/Q _6248_/A1 _5817_/A1 _7560_/Q _6333_/A1 _7800_/Q _4106_/A2 VDD VSS
+ gf180mcu_fd_sc_mcu7t5v0__aoi222_2
XFILLER_95_496 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_82_135 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7922_ _7922_/D _7923_/RN _7938_/CLK _7922_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
X_7853_ _7853_/D _7853_/RN _7853_/CLK _7853_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_82_179 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_36_574 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4996_ _3722_/I _3723_/I _5006_/B _5006_/C _4996_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__and4_4
X_7784_ _7784_/D _7901_/RN _7896_/CLK _7784_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffsnq_1
X_6804_ _7133_/S _6804_/A2 _6804_/B _7926_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_24_747 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6735_ _7761_/Q _6892_/A2 _6893_/C1 _7631_/Q _6738_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_3947_ _7788_/Q _6299_/A1 _5988_/A1 _7642_/Q _3948_/A4 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_149_432 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3878_ hold609/I _3869_/I _4231_/B1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_4
X_6666_ _7668_/Q _6891_/B1 _6880_/B1 _7806_/Q _6677_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_5617_ _5618_/B1 _5620_/B _5617_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__or2_1
X_6597_ _7912_/Q _7911_/Q _6953_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_4
X_5548_ _5548_/A1 _5548_/A2 _5548_/A3 _5765_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_136_159 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_151_129 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_145_682 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_144_170 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_132_321 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_117_384 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_3_629 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_5479_ _5779_/A1 _5479_/A2 _5503_/C VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_7218_ _7942_/Q _7228_/S _7219_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_120_527 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_7149_ _7699_/Q _7194_/A2 _7190_/B1 _7619_/Q _7153_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_86_463 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_58_176 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2135 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2113 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2124 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2102 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_104_85 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_104_96 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_104_74 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_64_34 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_61_308 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2168 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2157 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2146 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1423 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1412 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1401 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2179 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_154_2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1445 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1456 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1434 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1489 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1478 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1467 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_566 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_128_605 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_127_104 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_6_401 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_10_463 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_136_671 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_163_490 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_151_630 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_89_64 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_151_663 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_151_641 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_123_354 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_123_343 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_96_205 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_2_673 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_123_398 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_89_290 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_92_411 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_18_530 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_64_179 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_60_330 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4850_ hold47/Z _4852_/A2 _4850_/B _7509_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_45_382 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_159_730 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3801_ _3801_/I0 _3801_/I1 _3810_/S _3801_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_4
XFILLER_21_706 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1990 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_6520_ _6520_/A1 _6537_/A2 _6536_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_4
X_4781_ _6539_/A1 _4783_/A2 _4781_/B _7476_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_3732_ _7965_/Q _3731_/Z _3733_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_174_755 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_174_733 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_6451_ _6553_/A1 _6451_/A2 _6451_/B _7853_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_118_148 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3663_ _3663_/I _4392_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_9_283 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5402_ _5689_/A1 _5405_/B _5504_/A3 _5372_/Z _5576_/B2 _5577_/C VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai32_1
XFILLER_146_479 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_6382_ hold158/Z _6383_/A2 _6383_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_5333_ _5689_/A2 _5687_/B _5333_/A3 _5495_/B2 _5258_/B _5334_/C VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai32_1
XFILLER_127_682 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_114_321 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_114_343 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5264_ _5714_/B1 _5687_/B _5504_/A3 _5701_/C _5287_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai31_1
XFILLER_88_728 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5195_ _5087_/C _4914_/Z _5210_/A3 _5195_/B _5209_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai31_1
X_4215_ _7980_/Q _7965_/Q _7573_/Q _4215_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__or3_1
XFILLER_102_538 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7003_ _7003_/A1 _7133_/S _7003_/B1 _7003_/B2 _7932_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_68_463 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4146_ hold38/Z _4155_/A2 _4769_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_28_338 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_55_124 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4077_ input45/Z _4275_/A2 _5937_/A1 _7614_/Q _7646_/Q _6005_/A1 _4080_/A1 VDD VSS
+ gf180mcu_fd_sc_mcu7t5v0__aoi222_1
XFILLER_83_499 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_70_105 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7905_ _7905_/D _7961_/RN _7940_/CLK _7905_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_55_168 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_169_505 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_7836_ _7836_/D _7901_/RN _7854_/CLK _7836_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
Xclkbuf_leaf_96_csclk _7407_/CLK _7563_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_34_37 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_12_717 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4979_ _5069_/A2 _4930_/Z _4979_/A3 _4953_/Z _5366_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand4_4
XFILLER_11_227 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7767_ _7767_/D _7900_/RN _7767_/CLK _7767_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffsnq_1
X_7698_ _7698_/D _7853_/RN _7698_/CLK _7698_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
X_6718_ _7718_/Q _6881_/A2 _6885_/B1 _7710_/Q _6720_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_166_25 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_137_424 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_126_6 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6649_ _7910_/Q _6658_/A2 _6658_/A3 _6890_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor3_4
XFILLER_165_777 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_180_747 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xclkbuf_leaf_34_csclk clkbuf_3_7__f_csclk/Z _7726_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_133_641 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_160_460 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_59_89 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xclkbuf_leaf_49_csclk clkbuf_3_7__f_csclk/Z _7599_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_115_73 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_87_783 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_87_772 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_59_496 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_19_316 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_74_455 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_74_444 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_46_168 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_46_179 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_131_83 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1231 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1220 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_15_544 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_55_691 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1275 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1264 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1253 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1242 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1297 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1286 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_30_514 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_42_374 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_128_413 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xclkbuf_3_4__f_csclk clkbuf_0_csclk/Z _7873_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_30_569 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_156_744 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_11_783 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_6_231 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_109_682 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_171_769 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_170_246 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_136_490 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_111_302 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_97_503 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_85_709 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_69_238 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_111_357 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4000_ _4206_/A1 _7227_/I0 _4002_/B1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_93_753 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_92_241 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_65_499 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5951_ _4481_/I _5953_/A2 _5951_/B _7618_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_52_105 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4902_ _5309_/A1 _3723_/I _5666_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_5882_ hold770/Z _5885_/A2 _5883_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_7621_ _7621_/D _7961_/RN _7627_/CLK _7621_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffsnq_1
X_4833_ _6539_/A1 _4835_/A2 _4833_/B _7504_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_4764_ _4764_/A1 _6537_/A2 _4768_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_7552_ _7552_/D _7311_/Z _4418_/I1 _7552_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffnrnq_1
X_6503_ _6503_/A1 _6537_/A2 _6519_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_4
X_3715_ _7466_/Q _7184_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_7483_ _7483_/D _7949_/CLK _7483_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_4695_ hold617/Z _4718_/A1 _4698_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_119_479 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6434_ _6553_/A1 _6434_/A2 _6434_/B _7845_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_3646_ _7516_/Q _5678_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__inv_1
XFILLER_162_747 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_161_224 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_136_17 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_20_17 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_161_246 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6365_ hold313/Z _6366_/A2 _6366_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_115_641 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_142_460 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6296_ hold233/Z _6298_/A2 _6296_/B _7780_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_5316_ _5685_/B _5648_/B2 _5316_/B _5316_/C _5356_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi211_1
X_5247_ _5685_/B _5724_/B _5247_/B _5288_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
Xhold15 hold15/I hold15/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
Xhold37 hold37/I hold37/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
Xhold26 hold26/I hold26/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
X_5178_ _5178_/A1 _5178_/A2 _5178_/A3 _5188_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor3_1
Xhold59 hold59/I hold59/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
XFILLER_130_699 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_69_783 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xhold48 hold48/I hold48/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
XFILLER_28_124 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4129_ _4217_/A2 hold149/Z _4759_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_71_425 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_28_179 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_71_447 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_43_127 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_325 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_314 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_303 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_101_20 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_40_812 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_358 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_347 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_169_357 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_336 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
X_7819_ _7819_/D _7853_/RN _7821_/CLK _7819_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_61_35 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_138_755 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_20_580 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_137_298 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_137_276 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_117_2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_4_735 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_3_212 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_161_780 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_152_279 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_106_685 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_105_140 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_79_525 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_126_72 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_120_176 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_59_260 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_19_70 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_34_105 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_47_499 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_31_812 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_43_672 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_176_806 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1083 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1072 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1061 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1050 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_30_311 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_42_171 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_175_305 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1094 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_156_530 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_129_722 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_7_540 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4480_ hold232/Z hold49/Z _4480_/B hold233/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_4
XFILLER_167_90 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
Xhold507 hold507/I _4710_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
XFILLER_156_585 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_144_747 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xhold518 hold518/I _4498_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
XFILLER_7_562 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xhold529 _7602_/Q hold529/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
XFILLER_143_224 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_143_246 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_109_490 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6150_ hold600/Z _6157_/A2 hold601/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_98_812 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_801 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_5101_ _5602_/A1 _5647_/A2 _5777_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_2
XFILLER_32_2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_812 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_823 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_834 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_6081_ hold64/Z _6089_/A2 _6081_/B hold115/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
XTAP_845 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_856 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_867 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_5032_ _4965_/B _5366_/A2 _5608_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_4
XFILLER_111_176 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_78_591 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_878 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_889 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_57_219 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_81_712 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_65_274 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6983_ _7677_/Q _7191_/A2 _7191_/B1 _7799_/Q _6992_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_5934_ _4481_/I _5936_/A2 _5934_/B _7610_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_18_190 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_40_108 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_167_806 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5865_ hold637/Z _5868_/A2 _5866_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_22_812 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_179_699 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_178_176 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_178_165 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4816_ _4454_/Z _4816_/A2 _4816_/B _7495_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_7604_ _7604_/D _7961_/RN _7624_/CLK _7604_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffsnq_1
X_5796_ _5785_/B _5795_/Z _5806_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_4747_ _7460_/Q hold32/Z _4753_/S hold33/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_7535_ _7535_/D _7900_/RN _7823_/CLK _7535_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_162_522 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4678_ _7430_/Q _4685_/A1 _4681_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_7466_ _7466_/D _7900_/RN _7767_/CLK _7466_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
X_6417_ _6553_/A1 _6417_/A2 _6417_/B _7837_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_7397_ _7397_/D _7875_/RN _7823_/CLK _7397_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_122_408 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6348_ hold202/Z _6349_/A2 _6349_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_103_600 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_89_812 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_88_300 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_143_780 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xinput116 wb_adr_i[29] _4372_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyb_1
Xinput105 wb_adr_i[19] _4924_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyb_1
Xinput127 wb_cyc_i _4366_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XFILLER_130_463 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6279_ hold233/Z _6281_/A2 _6279_/B hold292/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_49_709 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xinput138 wb_dat_i[19] _7254_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyb_1
Xinput149 wb_dat_i[29] _7264_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XFILLER_56_46 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_57_753 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_57_764 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_16_105 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_29_477 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_72_756 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_29_499 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_112_63 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_72_34 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_100 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_71_288 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_133 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_122 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_13_812 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_111 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_169_176 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_166 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_155 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_144 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_12_333 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_199 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_188 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_177 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_172_308 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_153_544 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_126_747 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_141_739 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_141_706 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_137_60 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_106_460 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_98_108 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_97_97 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_153_70 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_121_496 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_63_712 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_90_531 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_35_425 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3980_ _7681_/Q _6073_/A1 hold28/I _7729_/Q _3981_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XPHY_2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_15_160 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_22_108 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5650_ _3728_/I _5122_/Z _5650_/A3 _5651_/A4 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_30_130 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_148_349 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4601_ _6539_/A1 _4603_/A2 _4601_/B _7403_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_5581_ _5212_/Z _5702_/A2 _5581_/B _5581_/C _5582_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XFILLER_129_563 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_7320_ _7877_/RN _4334_/Z _7320_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__and2_1
X_4532_ hold55/Z hold5/Z _4548_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_4
XFILLER_7_73 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_7251_ _7251_/A1 _7251_/A2 _7252_/C VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_4463_ hold49/Z _7258_/A1 _4464_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
Xhold315 _7731_/Q hold315/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
Xhold304 hold304/I _7715_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
Xhold326 _7673_/Q hold326/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
XFILLER_171_363 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_132_717 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
Xhold348 _7721_/Q hold348/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
XFILLER_117_19 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
Xhold337 hold337/I _7705_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
XFILLER_104_408 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6202_ _6547_/A1 _6208_/A2 _6202_/B hold556/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
Xhold359 hold359/I _7370_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
XFILLER_125_780 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4394_ _7444_/Q input80/Z _4396_/S _4394_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_7182_ _7182_/A1 _7182_/A2 _7182_/A3 _7183_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_97_152 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6133_ hold550/Z _6140_/A2 hold551/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_620 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_631 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_642 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_6064_ hold64/Z _6072_/A2 _6064_/B hold118/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_112_463 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_653 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_664 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_675 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_686 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_58_528 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5015_ _5139_/A1 _5014_/Z _5015_/B _5538_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi21_4
XTAP_697 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_38_230 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_81_531 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_38_274 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_53_211 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_54_723 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1819 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1808 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_26_469 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6966_ _7790_/Q _7190_/A2 _7194_/C1 _7806_/Q _6966_/C _6967_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi221_1
X_5917_ _4481_/I _5919_/A2 _5917_/B _7602_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_41_428 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_139_305 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6897_ _7210_/A1 _6767_/C _7433_/Q _6898_/B2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_179_496 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_139_316 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5848_ hold47/Z _5848_/A2 _5848_/B hold581/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_42_37 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_166_135 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_158_37 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5779_ _5779_/A1 _5779_/A2 _5779_/B1 _5292_/B _5780_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_7518_ _7518_/D _7959_/RN _7959_/CLK _7518_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_4
XFILLER_166_179 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_147_371 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_108_747 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_122_205 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_7449_ _7449_/D _7900_/RN _7887_/CLK _7449_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_174_69 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_162_396 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
Xhold860 _7740_/Q hold860/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
Xhold882 _7645_/Q hold882/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
Xhold871 _7783_/Q hold871/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
Xhold893 hold893/I _7526_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
XFILLER_131_783 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_130_282 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_103_496 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_67_89 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_29_230 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_123_40 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_76_369 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_29_241 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_45_712 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_123_73 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_83_22 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_17_425 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_44_200 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_45_778 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_60_737 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_157_113 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_13_686 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_8_123 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_172_105 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_141_503 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_126_577 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_114_717 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_99_428 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_4_362 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_79_141 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_95_601 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_35_211 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6820_ _7650_/Q _6880_/C2 _6892_/A2 _7764_/Q _6824_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_23_428 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6751_ hold79/I _6885_/A2 _6885_/B1 hold84/I _6752_/A4 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_3963_ _3783_/Z hold41/Z hold75/Z _3963_/A4 _3963_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__or4_2
XFILLER_16_480 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5702_ _5212_/Z _5702_/A2 _5702_/B _5702_/C _5782_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi211_2
X_3894_ _7805_/Q _6333_/A1 _5988_/A1 _7643_/Q _3896_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_6682_ _7798_/Q _6883_/A2 _6890_/B1 _7846_/Q _6683_/A4 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_148_157 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5633_ _5614_/Z _5622_/Z _5684_/A2 _5633_/A4 _5634_/A4 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand4_1
XFILLER_148_179 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5564_ _5565_/A1 _5565_/A2 _5565_/A3 _5578_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor3_1
Xhold101 _7817_/Q hold101/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
X_7303_ _7901_/RN _4334_/Z _7303_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__and2_1
X_4515_ _6547_/A1 _4521_/A2 _4515_/B hold651/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_160_812 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xhold112 hold112/I _7687_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
Xhold123 hold123/I _7695_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
X_5495_ _4993_/B _5647_/A2 _5797_/A2 _5687_/C _5495_/B2 _5742_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai32_1
Xhold134 _8005_/I hold134/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
X_7234_ _3658_/I _7281_/C2 _7235_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_4446_ hold49/I hold45/Z hold46/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
Xhold156 hold156/I _7723_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
Xhold167 _7841_/Q hold167/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
Xhold145 hold145/I _6511_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
X_4377_ _7965_/Q _4327_/S _4378_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_1
Xhold189 hold189/I _7691_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
Xhold178 hold178/I _7897_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
X_7165_ _7373_/Q _7203_/B1 _7204_/A2 _7399_/Q _7166_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_113_783 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_6116_ hold525/Z _6123_/A2 hold526/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_450 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_7096_ _7380_/Q _7188_/A2 _7096_/B _7097_/A4 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XTAP_494 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_483 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_461 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_472 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_6047_ hold64/Z _6055_/A2 _6047_/B _7663_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_100_477 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_85_144 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_27_712 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2317 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2306 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_54_531 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2339 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2328 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1605 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1649 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1638 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1627 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1616 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_7998_ _7998_/I _7998_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_6949_ _6949_/I _7210_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_3
XFILLER_10_601 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_167_499 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_154_105 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_127_308 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_10_656 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_6_605 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_154_127 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_108_544 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_151_812 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_123_503 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_108_566 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_108_555 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_78_33 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_162_193 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
Xhold690 _7578_/Q hold690/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
XFILLER_1_354 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_134_72 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_94_87 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_27_70 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_60_534 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_32_247 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_158_400 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_173_425 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_71_6 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_9_476 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
Xoutput217 _7991_/Z mgmt_gpio_out[17] VDD VSS gf180mcu_fd_sc_mcu7t5v0__buf_4
XFILLER_160_108 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_142_812 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xoutput206 _3705_/ZN mgmt_gpio_oeb[7] VDD VSS gf180mcu_fd_sc_mcu7t5v0__buf_4
XFILLER_57_4 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4300_ _3812_/Z _4297_/Z _4300_/B _4300_/C _4301_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai211_1
Xoutput239 _4386_/Z mgmt_gpio_out[37] VDD VSS gf180mcu_fd_sc_mcu7t5v0__buf_4
Xoutput228 _8001_/Z mgmt_gpio_out[27] VDD VSS gf180mcu_fd_sc_mcu7t5v0__buf_4
XFILLER_126_396 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_114_514 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5280_ _5482_/B2 _5292_/B _5690_/A1 _5575_/A2 _5412_/B _5282_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi221_1
XFILLER_5_682 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_4231_ input71/Z _5903_/A1 _4231_/B1 input36/Z _4280_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_141_377 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_141_366 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_4_63 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4162_ _4162_/A1 _4162_/A2 _4162_/A3 _4204_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand3_1
X_4093_ _7816_/Q _6367_/A1 _6316_/A1 _7792_/Q _5870_/A1 _7577_/Q _4106_/A1 VDD VSS
+ gf180mcu_fd_sc_mcu7t5v0__aoi222_2
XFILLER_67_144 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_28_509 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_7921_ _7921_/D _7938_/RN _7938_/CLK _7921_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_36_531 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7852_ _7852_/D _7877_/RN _7852_/CLK _7852_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_51_512 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_51_523 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_4995_ _5602_/A2 _4993_/B _4993_/C _4998_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor3_1
XFILLER_91_692 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_90_191 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6803_ _7926_/Q _7133_/S _6804_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_63_383 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7783_ _7783_/D _7900_/RN _7900_/CLK _7783_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffsnq_1
X_6734_ hold69/I _6892_/B1 _6738_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_3946_ _7618_/Q _5937_/A1 _6226_/A1 _7754_/Q _7804_/Q _6333_/A1 _3948_/A3 VDD VSS
+ gf180mcu_fd_sc_mcu7t5v0__aoi222_2
XFILLER_51_567 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_177_753 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_139_39 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_136_105 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3877_ hold38/Z _3847_/Z _6005_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_4
X_6665_ _7910_/Q _6665_/A2 _6665_/A3 _6665_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__and3_2
XFILLER_149_499 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5616_ _5616_/A1 _5643_/B1 _5176_/B _5620_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor3_4
X_6596_ _7434_/Q _6599_/A2 _6596_/B _7911_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_5547_ _5547_/A1 _5547_/A2 _5764_/A2 _5646_/A2 _5549_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor4_1
XFILLER_133_812 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5478_ _5797_/A1 _5543_/C _5543_/B _5545_/B _5662_/A1 _5505_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai32_1
XFILLER_105_514 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_144_193 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7217_ _7517_/D _7959_/RN _7228_/S VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_4
X_4429_ _4400_/S input68/Z _4429_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__and2_1
X_7148_ _7148_/A1 _7148_/A2 _7148_/A3 _7159_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_101_753 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_7079_ _7079_/A1 _7210_/A2 _7433_/Q _7080_/B2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XTAP_2114 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2125 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2103 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2158 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2147 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2136 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1424 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1413 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1402 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_64_46 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_15_704 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_54_372 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_2169 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1446 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1457 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1435 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_14_247 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_42_534 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_147_2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1479 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1468 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_168_742 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_80_56 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_22_291 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_155_436 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_155_425 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_182_244 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_142_108 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_129_83 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_135_160 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_124_812 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_89_54 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_89_87 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_89_280 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_49_144 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_49_199 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_18_542 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_52_309 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_18_597 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3800_ hold49/Z _3801_/I1 _3800_/B hold53/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_4
X_4780_ hold738/Z _4783_/A2 _4781_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_33_567 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1991 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1980 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_3731_ _3744_/A1 _7411_/Q _3730_/Z _3731_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__and3_1
XFILLER_158_252 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xclkbuf_leaf_0_csclk _7407_/CLK _7823_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
X_3662_ _3662_/I _4380_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_6450_ hold314/Z _6451_/A2 _6451_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_118_116 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5401_ _5673_/A1 _5706_/A2 _5401_/A3 _5401_/A4 _5414_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand4_1
XFILLER_62_2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6381_ _4481_/I _6383_/A2 _6381_/B _7820_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_161_428 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_115_812 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_114_311 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_5332_ _5258_/B _5495_/B2 _5757_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_130_804 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_114_333 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_5_490 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_125_19 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5263_ _5433_/C _5768_/A3 _5681_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_5194_ _5199_/B _3727_/I _4915_/Z _4996_/Z _5371_/C VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand4_4
X_4214_ _3828_/I _4075_/B _5852_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_87_228 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7002_ _7931_/Q _6556_/B _7002_/B _7003_/B2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_4145_ hold38/Z _3869_/I _4843_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_95_283 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_95_272 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_83_412 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_83_423 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4076_ _7880_/Q _6503_/A1 _4104_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_7904_ _7904_/D _7961_/RN _7940_/CLK _7904_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
X_7835_ _7835_/D _7901_/RN _7901_/CLK _7835_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_70_128 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_24_534 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_36_383 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4978_ _5104_/B _5669_/B _4999_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_7766_ _7766_/D _7900_/RN _7767_/CLK _7766_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffsnq_1
XFILLER_51_397 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_165_712 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_7697_ _7697_/D _7923_/RN _7698_/CLK _7697_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
X_6717_ _7646_/Q _6880_/C2 _6882_/B1 _7654_/Q _6720_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_3929_ hold76/I _4075_/B _4176_/C VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_164_211 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_20_784 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6648_ _6878_/A2 _6663_/A4 _6664_/A2 _6880_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor3_4
XFILLER_50_37 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_166_37 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_165_767 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_164_266 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_137_469 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_124_119 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_124_108 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_117_160 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6579_ _7907_/Q _7906_/Q _6663_/A4 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_4
XFILLER_182_69 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_182_47 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_78_239 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_59_79 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_86_250 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_115_96 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_47_648 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_46_125 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_131_73 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_1232 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1221 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1210 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_61_139 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_91_66 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_91_44 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_1265 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1254 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1243 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_70_673 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_15_567 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_42_364 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1298 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1287 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1276 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_70_695 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_128_403 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_156_756 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_11_762 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_10_250 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_128_458 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_116_609 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_6_243 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_143_428 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_123_141 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_123_174 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_69_228 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_2_460 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_2_471 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_78_795 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_77_283 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_65_423 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_93_776 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5950_ hold708/Z _5953_/A2 _5951_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_4901_ _3722_/I _5006_/B _5006_/C _4946_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand3_4
XFILLER_80_459 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_61_651 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7620_ _7620_/D _7961_/RN _7624_/CLK _7620_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffsnq_1
X_5881_ _5881_/A1 _6537_/A2 _5885_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_4832_ hold755/Z _4835_/A2 _4833_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_159_550 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_147_712 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4763_ _4454_/Z _4763_/A2 _4763_/B _7469_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_7551_ _7551_/D _7310_/Z _4418_/I1 _7551_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffnrnq_1
XFILLER_174_531 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_146_211 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6502_ _6553_/A1 _6502_/A2 _6502_/B hold311/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_4694_ _4718_/A1 _4694_/A2 _4694_/B hold616/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_119_425 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3714_ _7611_/Q _6849_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_7482_ _7482_/D _7949_/CLK _7482_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_6433_ hold250/Z _6434_/A2 _6434_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_174_575 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3645_ _7517_/Q _4376_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_106_108 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_6364_ hold233/Z _6366_/A2 _6364_/B _7812_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_6295_ hold389/Z _6298_/A2 _6296_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_5315_ _5545_/A2 _5687_/B _5648_/B2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_4
XFILLER_0_419 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5246_ _5199_/B _5201_/B _5421_/A1 _5333_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand3_1
Xhold16 hold16/I hold16/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
Xhold27 hold27/I hold27/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
Xhold38 hold38/I hold38/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
XFILLER_102_369 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_69_773 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
Xhold49 hold49/I hold49/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
X_5177_ _5651_/A1 _5769_/A1 _5177_/A3 _5178_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_68_250 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_29_637 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_29_626 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4128_ _4141_/A1 _4151_/A2 _4868_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_4059_ _7849_/Q _6435_/A1 _6265_/A1 _7769_/Q _4232_/A2 input6/Z _4063_/A1 VDD VSS
+ gf180mcu_fd_sc_mcu7t5v0__aoi222_1
XFILLER_83_286 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_315 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_304 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_101_43 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XPHY_359 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_348 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_337 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_326 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_101_65 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_7818_ _7818_/D _7853_/RN _7818_/CLK _7818_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_24_375 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_51_150 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_52_673 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_52_684 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7749_ _7749_/D _7877_/RN _7809_/CLK _7749_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffsnq_1
XFILLER_138_723 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_138_767 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_165_586 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_125_428 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_180_534 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_152_247 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_4_747 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_126_84 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_86_33 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_86_44 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_87_570 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_47_423 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_75_743 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_59_283 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_142_72 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_47_478 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_90_735 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_34_117 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_1040 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_15_353 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_35_70 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1073 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1062 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1051 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_129_712 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_70_492 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1095 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1084 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_128_211 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_30_389 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xclkbuf_leaf_80_csclk clkbuf_leaf_9_csclk/I _7847_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_11_570 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xhold508 hold508/I _7441_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
Xhold519 hold519/I _7359_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
XFILLER_171_578 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_171_567 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xclkbuf_leaf_95_csclk _7407_/CLK _7567_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
X_6080_ hold113/Z _6089_/A2 hold114/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_5100_ _5705_/A2 _5585_/A1 _5573_/C _5105_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XTAP_802 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_813 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_824 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_835 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_111_144 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_5031_ _5104_/B _5658_/B _5031_/B _5038_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_85_507 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_846 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_857 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_868 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_25_2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_879 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_65_286 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_25_139 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6982_ _7791_/Q _7190_/A2 _7190_/B1 _7613_/Q _7190_/C1 _7701_/Q _6992_/A2 VDD VSS
+ gf180mcu_fd_sc_mcu7t5v0__aoi222_1
Xclkbuf_leaf_33_csclk clkbuf_3_7__f_csclk/Z _7811_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
X_5933_ hold711/Z _5936_/A2 _5934_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_5864_ _6549_/A1 _5868_/A2 _5864_/B _7578_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_34_673 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_179_689 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_7603_ hold10/Z _7853_/RN _7603_/CLK hold8/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
X_4815_ hold813/Z _4816_/A2 _4816_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_5795_ _5795_/A1 _5795_/A2 _5795_/A3 _5795_/A4 _5795_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__or4_1
X_7534_ _7534_/D _7961_/RN _7650_/CLK _7534_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
Xclkbuf_leaf_48_csclk clkbuf_3_7__f_csclk/Z _7603_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_147_564 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4746_ _4454_/Z _4753_/S _4746_/B _7459_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_7465_ _7465_/D _7853_/RN _7601_/CLK _7465_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
X_4677_ _4685_/A1 _4677_/A2 _4677_/B hold613/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_107_428 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_162_534 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_134_247 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6416_ hold246/Z _6417_/A2 _6417_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_7396_ _7396_/D _7961_/RN _7401_/CLK _7396_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
X_6347_ hold233/Z _6349_/A2 _6347_/B _7804_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_88_323 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xinput117 wb_adr_i[2] _5006_/C VDD VSS gf180mcu_fd_sc_mcu7t5v0__buf_12
Xinput106 wb_adr_i[1] _3722_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__buf_12
XFILLER_103_645 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_88_367 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6278_ hold291/Z _6281_/A2 _6279_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
Xinput128 wb_dat_i[0] _7242_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyb_1
Xinput139 wb_dat_i[1] _7247_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XFILLER_102_188 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5229_ _5290_/B _5645_/A3 _5573_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_88_389 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_69_570 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_17_618 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_112_31 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_71_223 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_71_212 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_44_426 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_134 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_123 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_101 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_112 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_169_144 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_167 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_156 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_145 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_24_183 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_189 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_178 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_40_676 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_138_531 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_12_389 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_125_236 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_180_353 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_153_567 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_141_718 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_79_312 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_94_315 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_772 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_35_415 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_47_286 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_62_245 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_35_448 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_35_459 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_16_673 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_149_807 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4600_ hold766/Z _4603_/A2 _4601_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_5580_ _5580_/A1 _5636_/A1 _5380_/I _5581_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__or3_1
X_4531_ _4454_/Z _4531_/A2 _4531_/B _7374_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_7250_ _7520_/Q _7250_/A2 _7250_/B1 _7518_/Q _7251_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_144_534 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
Xhold316 _7797_/Q hold316/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
Xhold305 _7836_/Q hold305/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
X_4462_ _4487_/A1 _4460_/Z _4462_/B _7349_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
Xhold327 hold327/I _6068_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
Xhold338 _7745_/Q hold338/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
Xhold349 hold349/I _7721_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
XFILLER_116_258 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_116_247 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_89_109 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6201_ hold554/Z _6208_/A2 hold555/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_125_792 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_4393_ _7881_/Q _4396_/S _4393_/B _4393_/ZN VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_7181_ _7371_/Q _7201_/A2 _7205_/B1 _7537_/Q _7182_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_6132_ hold64/Z _6140_/A2 _6132_/B hold126/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_98_676 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_610 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_621 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_632 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_643 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_6063_ hold116/Z _6072_/A2 hold117/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_100_626 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_100_615 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_97_164 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_654 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_665 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_676 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_5014_ _5195_/B _4926_/Z _5010_/Z _5014_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__or3_2
XTAP_687 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_698 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_38_220 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_93_392 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_26_28 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_26_17 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1809 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_26_448 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6965_ _6965_/A1 _6965_/A2 _6965_/A3 _6966_/C VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand3_1
X_5916_ hold529/Z _5919_/A2 _5917_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_81_587 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_41_418 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_21_120 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_6896_ _6888_/Z _6896_/A2 _6896_/A3 _6895_/Z _6898_/B1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand4_1
X_5847_ _7571_/Q _5848_/A2 _5848_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_22_676 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5778_ _5778_/A1 _5737_/B _5710_/Z _5733_/Z _5785_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__and4_1
XFILLER_21_175 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_21_164 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_182_629 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7517_ _7517_/D _7959_/RN _7959_/CLK _7517_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_163_810 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_147_361 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4729_ _6547_/A1 _4731_/A2 _4729_/B hold457/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_108_737 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_107_225 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_7448_ _7448_/D _7900_/RN _7887_/CLK _7448_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_174_37 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_135_567 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_123_707 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7379_ hold56/Z _7877_/RN _7381_/CLK _7379_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_1_525 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
Xhold861 _7394_/Q hold861/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
Xhold850 _7536_/Q hold850/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
Xhold872 _7839_/Q hold872/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
Xhold894 _7629_/Q hold894/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
Xhold883 _7605_/Q hold883/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
XFILLER_130_250 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_49_507 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_49_518 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_177_2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_83_34 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_29_286 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_44_212 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_84_392 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_44_256 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_72_576 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_60_727 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_9_636 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_8_135 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_40_495 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_8_179 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_32_60 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_166_692 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_148_82 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_126_534 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_126_523 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_121_283 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_83_808 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_82_318 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_94_189 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_75_392 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_36_757 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6750_ hold66/I _6644_/Z _6884_/B1 _7687_/Q _6752_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_5701_ _5405_/B _5701_/A2 _5780_/A2 _5382_/Z _5701_/C _5702_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai221_2
XFILLER_92_2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3962_ input31/Z _4249_/A2 _5870_/A1 _3961_/Z _3998_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_148_114 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3893_ _7667_/Q _6039_/A1 _6022_/A1 _7659_/Q _6056_/A1 _7675_/Q _3896_/A1 VDD VSS
+ gf180mcu_fd_sc_mcu7t5v0__aoi222_2
X_6681_ _6681_/A1 _6681_/A2 _6681_/A3 _6681_/A4 _6684_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand4_1
X_5632_ _5632_/A1 _5632_/A2 _5697_/A2 _5697_/A3 _5633_/A4 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor4_1
XFILLER_163_106 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_145_810 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5563_ _5663_/A1 _5405_/B _5381_/Z _5618_/B1 _5563_/B2 _5565_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai32_1
XFILLER_117_501 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_12_19 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_7302_ _7901_/RN _4334_/Z _7302_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__and2_1
X_4514_ hold649/Z _4521_/A2 hold650/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_5494_ _5648_/A1 _5658_/B _5176_/B _5425_/B _5767_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_1
Xhold124 _7703_/Q hold124/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
XFILLER_117_567 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xhold113 _7679_/Q hold113/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
XFILLER_105_707 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
Xhold102 _7785_/Q hold102/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
Xhold135 hold135/I _5902_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
X_7233_ _7520_/Q _7233_/A2 _7233_/B1 _7518_/Q _7238_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_2
Xhold168 _7777_/Q hold168/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
X_4445_ hold840/Z _4487_/A1 _4450_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
Xhold157 _7561_/Q hold157/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
Xhold146 hold146/I _7881_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
X_4376_ _7214_/A1 _7214_/A2 _4376_/B _7511_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
Xhold179 _7639_/Q hold179/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
X_7164_ _7403_/Q _7203_/A2 _7204_/B1 _7389_/Q _7166_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_112_250 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_6115_ hold64/Z _6123_/A2 _6115_/B hold123/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_98_473 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_98_484 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_86_624 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_86_602 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_451 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_440 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_98_495 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7095_ _7095_/A1 _7095_/A2 _7096_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_484 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_462 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_473 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_6046_ hold79/Z _6055_/A2 _6047_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_100_467 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_495 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2307 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_54_521 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2329 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2318 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1606 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_66_392 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7997_ _7997_/I _7997_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_1639 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1628 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1617 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_41_215 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6948_ _6955_/A4 _6948_/A2 _6946_/Z _6948_/A4 _6949_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand4_4
XFILLER_22_451 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6879_ _6879_/A1 _6879_/A2 _6889_/C VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_139_136 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_10_646 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_108_534 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_2_812 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_150_334 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
Xhold680 hold680/I _6109_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
XFILLER_150_389 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_131_570 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_1_366 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
Xhold691 _7652_/Q hold691/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
XFILLER_103_294 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_103_283 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_76_134 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_92_605 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_77_668 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_65_808 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_92_627 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_64_318 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_17_212 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_45_532 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_57_392 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_60_524 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_60_579 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_60_568 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_32_259 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_43_70 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_159_70 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_139_692 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_9_499 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xoutput207 _3704_/ZN mgmt_gpio_oeb[8] VDD VSS gf180mcu_fd_sc_mcu7t5v0__buf_4
Xoutput218 _7992_/Z mgmt_gpio_out[18] VDD VSS gf180mcu_fd_sc_mcu7t5v0__buf_4
XFILLER_154_673 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xoutput229 _8002_/Z mgmt_gpio_out[28] VDD VSS gf180mcu_fd_sc_mcu7t5v0__buf_4
XFILLER_99_215 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_114_548 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4230_ _7546_/Q _5807_/A1 _5871_/A1 _7582_/Q _4280_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_68_602 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4161_ _7669_/Q _6056_/A1 _4764_/A1 _7471_/Q _4162_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_4092_ _4084_/Z _4092_/A2 _4092_/A3 _4092_/A4 _4107_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand4_2
XFILLER_83_638 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7920_ _7920_/D _7961_/RN _7940_/CLK _7920_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
X_7851_ _7851_/D _7853_/RN _7851_/CLK _7851_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_48_392 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6802_ _7433_/Q _7925_/Q _6802_/B1 _6802_/B2 _6804_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_91_682 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4994_ _5602_/A2 _4993_/B _5648_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_2
XFILLER_90_181 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_23_215 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7782_ _7782_/D _7900_/RN _7900_/CLK _7782_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffsnq_1
X_6733_ _7133_/S _6733_/A2 _6733_/B _7923_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_3945_ input50/Z _4275_/A2 _4231_/B1 input69/Z _3948_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_6664_ _6878_/A2 _6664_/A2 _6664_/A3 _6880_/B1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor3_4
X_5615_ _5689_/A1 _5692_/B _5618_/A3 _5763_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor3_2
X_3876_ hold72/Z hold38/Z _5971_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_4
XFILLER_31_292 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_136_139 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_6595_ _6599_/A2 _6618_/A3 _6596_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_164_459 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5546_ _5797_/A2 _5546_/A2 _5546_/B1 _5543_/B _5546_/C _5646_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai221_2
XFILLER_133_802 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_160_621 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_144_150 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5477_ _5496_/A1 _5797_/B _4965_/B _5543_/B _5477_/B2 _5510_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai32_1
XFILLER_2_108 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7216_ _7216_/A1 _7216_/A2 _7941_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_4428_ _4428_/I _7963_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_160_676 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xclkbuf_2_3__f_mgmt_gpio_in[4] clkbuf_0_mgmt_gpio_in[4]/Z _7972_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_132_389 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_59_602 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_113_570 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7147_ _7683_/Q _7191_/A2 _6938_/I _7861_/Q _7148_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_4359_ _4361_/A3 _4359_/A2 _4359_/B _7434_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_48_37 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_104_21 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_86_465 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7078_ _7210_/A2 _7078_/A2 _7078_/A3 _7078_/A4 _7078_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__or4_1
XFILLER_74_605 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_47_808 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_58_134 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6029_ hold127/Z _6038_/A2 _6030_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_46_318 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2115 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2126 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2104 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_39_392 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_2159 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2148 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2137 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1414 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1403 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_70_800 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_1447 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1436 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1425 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_120_42 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_1469 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1458 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_14_259 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_128_607 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_80_68 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_182_212 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_167_286 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_13_73 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_129_73 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_129_62 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_6_458 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_182_278 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_136_673 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_123_301 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_1_141 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_2_664 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_145_83 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_89_292 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_77_465 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_77_454 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_77_443 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_38_808 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_77_487 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_65_638 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_61_811 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_60_321 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_60_310 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_45_384 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_178_529 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1970 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_3730_ _7346_/Q _7345_/Q _3730_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__and2_1
XTAP_1992 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1981 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_173_212 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3661_ _3661_/I _4368_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_5400_ _5585_/A1 _5658_/B _5685_/B _5759_/A1 _5401_/A4 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_6380_ hold715/Z _6383_/A2 _6381_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_9_296 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5331_ _5645_/A1 _5687_/B _5618_/A3 _5331_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__or3_1
XFILLER_55_2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_142_676 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_5262_ _5687_/B _5504_/A3 _5779_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_7001_ _7605_/Q _6949_/I _7001_/B1 _7001_/B2 _7001_/C _7003_/B1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai221_1
X_5193_ _5199_/B _4915_/Z _4996_/Z _5202_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_114_389 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4213_ _7652_/Q _6022_/A1 _4843_/A1 _7507_/Q _4262_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_4144_ input44/Z _4275_/A2 _4719_/A1 input62/Z _4198_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_29_808 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_56_605 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_110_584 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_28_318 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4075_ hold76/I _3963_/Z _4075_/B _4083_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_7903_ _7903_/D _7961_/RN _7940_/CLK _7903_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
X_7834_ _7834_/D _7901_/RN _7878_/CLK _7834_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_63_170 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_34_17 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7765_ _7765_/D _7853_/RN _7851_/CLK _7765_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_51_354 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_177_540 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4977_ _5603_/A1 _4993_/B _5669_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_4
X_6716_ _6716_/A1 _6716_/A2 _6716_/A3 _6716_/A4 _6721_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand4_1
XFILLER_11_229 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3666__1 _3666__1/I _7279_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_7696_ _7696_/D _7923_/RN _7720_/CLK _7696_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
X_3928_ _7796_/Q _6316_/A1 _3943_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_164_201 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_149_286 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_109_106 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3859_ hold89/Z _4141_/A1 hold90/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_4
X_6647_ _6878_/A2 _6665_/A2 _6665_/A3 _6647_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__and3_2
XFILLER_164_256 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6578_ _4352_/B _7907_/Q _6581_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_5529_ _5201_/B _5529_/A2 _5529_/A3 _5548_/A3 _5541_/A4 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand4_2
XFILLER_118_673 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_117_172 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_3_428 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_182_37 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_132_197 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_132_186 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_86_273 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_74_402 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_75_24 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_59_476 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_19_307 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_47_638 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1222 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1211 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1200 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_321 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_131_96 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_91_56 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1266 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1255 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1244 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1233 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1299 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1288 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1277 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_24_61 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_156_735 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_155_223 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_155_212 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_7_712 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_143_407 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_115_109 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_6_277 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_170_259 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_124_676 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_38_605 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_1_32 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_93_799 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_65_479 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4900_ _3722_/I _5006_/B _5006_/C _4900_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__and3_2
X_5880_ hold47/Z _5880_/A2 _5880_/B _7585_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_65_90 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_46_693 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_61_641 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4831_ _4831_/A1 _6537_/A2 _4835_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_33_354 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_33_343 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_159_540 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_147_702 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_4762_ hold889/Z _4763_/A2 _4763_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_7550_ _7550_/D _7309_/Z _4418_/I1 _7550_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffnrnq_1
XFILLER_174_521 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6501_ hold309/Z _6502_/A2 hold310/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_4693_ hold615/Z _3819_/Z _4693_/B _4694_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_3713_ _7610_/Q _6826_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_7481_ _7481_/D _7949_/CLK _7481_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_3644_ _7411_/Q _4292_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__inv_3
X_6432_ hold233/Z _6434_/A2 _6432_/B hold284/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_161_215 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_161_248 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6363_ hold390/Z _6366_/A2 _6364_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_130_602 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6294_ _6549_/A1 _6298_/A2 _6294_/B _7779_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_5314_ _5692_/B _5365_/B1 _5618_/A3 _5316_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor3_1
X_5245_ _3728_/I _5369_/B _5271_/A3 _5724_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor3_4
XFILLER_69_730 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
Xhold17 hold17/I hold17/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
Xhold28 hold28/I hold28/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
XFILLER_130_646 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_114_197 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5176_ _5027_/Z _5479_/A2 _5176_/B _5177_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
Xhold39 hold39/I hold39/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
XFILLER_110_392 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_84_744 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_84_733 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_83_232 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4127_ _7749_/Q _6226_/A1 _4158_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_4058_ _4058_/A1 _4058_/A2 _4058_/A3 _4058_/A4 _4069_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor4_2
XFILLER_84_788 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_71_405 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_316 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_305 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_24_321 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_349 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_338 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_327 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
X_7817_ _7817_/D _7853_/RN _7821_/CLK _7817_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_24_387 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_52_696 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_7748_ _7748_/D _7877_/RN _7755_/CLK _7748_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffsnq_1
XFILLER_137_212 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_131_6 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7679_ _7679_/D _7923_/RN _7735_/CLK _7679_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_137_223 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_153_738 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_3_225 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_106_676 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_105_164 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_120_123 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_86_23 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_120_189 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_19_104 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_101_392 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_74_265 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_16_800 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_90_747 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_62_449 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_27_170 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1030 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_43_641 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_70_471 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_70_460 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1074 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1063 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1052 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1041 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_30_302 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1096 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1085 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_175_318 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_168_392 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_51_70 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_167_70 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_116_407 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
Xhold509 _7658_/Q hold509/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
XFILLER_171_557 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_143_248 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_143_215 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_152_771 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_112_602 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_803 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_814 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_825 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_5030_ _5496_/A1 _5458_/C _5661_/A1 _5031_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor3_1
XFILLER_97_357 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_836 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_847 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_858 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_869 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_66_744 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_18_2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_38_424 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_66_788 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6981_ _7709_/Q _7189_/A2 _7189_/B1 _7685_/Q _7189_/C1 _7653_/Q _6992_/A1 VDD VSS
+ gf180mcu_fd_sc_mcu7t5v0__aoi222_1
X_5932_ _4476_/I _5936_/A2 _5932_/B hold342/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_19_682 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_15_19 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_18_181 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_18_192 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5863_ hold690/Z _5868_/A2 _5864_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_21_302 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_178_145 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7602_ _7602_/D _7853_/RN _7603_/CLK _7602_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
X_5794_ _5794_/A1 _5794_/A2 _5794_/A3 _5795_/A4 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand3_1
X_4814_ hold47/Z _4816_/A2 _4814_/B hold411/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_33_195 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_166_318 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4745_ hold618/Z _4753_/S _4746_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_119_212 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_21_357 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7533_ _7533_/D _7961_/RN _7572_/CLK _7533_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
X_7464_ _7464_/D _7853_/RN _7601_/CLK _7464_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
X_4676_ _7463_/Q _3879_/Z _4676_/B _4677_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_6415_ hold233/Z _6417_/A2 _6415_/B hold306/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_7395_ _7395_/D _7938_/RN _7401_/CLK _7395_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
X_6346_ hold371/Z _6349_/A2 _6347_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_142_270 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_115_495 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_228 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
Xinput107 wb_adr_i[20] _5195_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_8
Xinput118 wb_adr_i[30] _4367_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyb_1
X_6277_ _6549_/A1 _6281_/A2 _6277_/B _7771_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
Xinput129 wb_dat_i[10] _7249_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyb_1
X_5228_ _5200_/B _3727_/I _3728_/I _5022_/B _5645_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand4_4
XFILLER_130_487 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5159_ _4965_/B _5366_/A2 _5797_/A2 _5752_/C VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor3_2
XFILLER_56_37 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_56_59 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_57_777 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_72_747 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_72_736 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_25_641 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_169_101 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_124 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_24_162 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_102 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_52_460 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_113 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_157 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_146 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_135 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_179 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_168 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_8_317 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_138_543 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_138_521 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_122_2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_181_800 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_138_587 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_180_321 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_137_40 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_125_215 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_4_534 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_21_73 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_137_73 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_137_51 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_134_760 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_137_95 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_106_484 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_106_473 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_106_495 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_97_99 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_97_77 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_95_806 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_79_357 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_121_454 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_153_83 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_48_744 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_48_766 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_90_544 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_63_769 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_71_780 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_4 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_43_460 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_50_419 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_176_605 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_148_329 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_148_318 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_169_690 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_30_176 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_31_699 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4530_ hold863/Z _4531_/A2 _4531_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_4461_ _4461_/A1 hold31/Z hold32/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
Xhold317 hold317/I _6332_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
Xhold306 hold306/I _7836_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
XFILLER_171_354 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xhold339 hold339/I _7745_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
Xhold328 hold328/I _7673_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
X_6200_ hold64/Z _6208_/A2 _6200_/B hold130/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_7180_ _7960_/Q _7207_/A2 _7207_/B1 _7529_/Q _7205_/A2 _7533_/Q _7182_/A2 VDD VSS
+ gf180mcu_fd_sc_mcu7t5v0__aoi222_1
X_6131_ hold124/Z _6140_/A2 hold125/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_600 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_4392_ _4392_/A1 _4396_/S _4393_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_140_741 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_611 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_622 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_633 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_100_605 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_97_176 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6062_ _4460_/Z _6072_/A2 _6062_/B _7670_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
XTAP_644 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_655 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_666 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_677 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_5013_ _5195_/B _4926_/Z _5010_/Z _5016_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor3_2
XFILLER_112_498 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_85_327 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_688 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_699 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_39_722 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_66_585 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_39_799 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_54_747 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6964_ _7878_/Q _7203_/B1 _7193_/C1 _7724_/Q _6965_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_5915_ _4476_/I _5919_/A2 _5915_/B hold221/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_34_460 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6895_ _6895_/A1 _6895_/A2 _6895_/A3 _6895_/A4 _6895_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__and4_1
XFILLER_179_454 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5846_ hold580/Z _7285_/A2 _5848_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_42_17 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_139_307 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5777_ _5777_/A1 _5777_/A2 _5777_/B _5777_/C _5802_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi211_2
X_7516_ _7516_/D _7959_/RN _7959_/CLK _7516_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
X_4728_ hold455/Z _4731_/A2 hold456/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_175_682 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_162_321 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4659_ _3879_/Z _4454_/Z _4660_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_107_215 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_7447_ _7447_/D _7875_/RN _7881_/CLK _7447_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
X_7378_ _7378_/D _7877_/RN _7752_/CLK _7378_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_162_398 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_162_376 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
Xhold840 _7347_/Q hold840/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
Xhold862 _7587_/Q hold862/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
Xhold851 _7392_/Q hold851/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
Xhold873 _7831_/Q hold873/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
Xhold895 _7376_/Q hold895/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
XFILLER_89_655 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6329_ hold710/Z _6332_/A2 _6330_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
Xhold884 _7637_/Q hold884/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
XFILLER_88_176 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_88_198 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_29_221 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_29_232 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_123_86 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_123_97 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_60_717 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_158_605 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_13_611 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
Xclkbuf_leaf_94_csclk _7407_/CLK _7875_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_53_780 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_40_463 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_157_126 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_12_176 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_138_351 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_181_641 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_180_140 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_153_354 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xclkbuf_leaf_32_csclk clkbuf_3_6__f_csclk/Z _7805_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_106_270 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_164_71 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_95_603 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_121_295 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_94_124 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_94_102 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xclkbuf_leaf_47_csclk clkbuf_3_7__f_csclk/Z _7419_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_36_703 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_94_179 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_36_747 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_63_577 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3961_ _7930_/Q _7578_/Q _7580_/Q _3961_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_16_460 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_35_279 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5700_ _5104_/B _5212_/Z _5780_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_16_471 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_149_638 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_148_104 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3892_ _3892_/A1 _3892_/A2 _3892_/A3 _3892_/A4 _3918_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand4_2
X_6680_ _7716_/Q _6881_/A2 _6885_/A2 _7660_/Q _6681_/A4 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_5631_ _5331_/Z _5437_/B _5619_/Z _5697_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_85_2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_31_496 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5562_ _5735_/A2 _5585_/A1 _5562_/B _5704_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_7301_ _7901_/RN _4334_/Z _7301_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_144_321 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4513_ _6545_/A1 _4521_/A2 _4513_/B hold287/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_7232_ _3658_/I _7281_/B1 _7233_/B1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
Xhold114 hold114/I _6081_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
X_5493_ _5603_/A1 _4993_/B _5797_/A2 _5493_/B _5530_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai31_1
Xhold125 hold125/I _6132_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
Xhold103 hold103/I _7785_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
Xhold147 _7340_/Q hold147/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
Xhold158 _7821_/Q hold158/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
Xhold136 hold136/I _7595_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
X_4444_ hold194/Z _6537_/A2 _4487_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_4
X_4375_ _4375_/A1 _4375_/A2 _7214_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_144_19 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
Xhold169 _7801_/Q hold169/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
X_7163_ _7407_/Q _7202_/A2 _7202_/B1 _7397_/Q _7385_/Q _7202_/C2 _7166_/A1 VDD VSS
+ gf180mcu_fd_sc_mcu7t5v0__aoi222_1
X_6114_ hold121/Z _6123_/A2 hold122/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_98_463 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7094_ _7899_/Q _7197_/A2 _6938_/I _7859_/Q _7095_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XTAP_441 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_430 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_6045_ _4460_/Z _6055_/A2 _6045_/B _7662_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
XTAP_485 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_463 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_474 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_452 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_85_168 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_496 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_37_17 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2308 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_26_202 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_39_574 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2319 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_26_246 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_27_769 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_54_544 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_7996_ _7996_/I _7996_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_1629 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1618 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1607 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_54_566 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6947_ _7195_/A2 _7195_/C1 _7207_/B1 _7196_/B1 _6948_/A4 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor4_4
XFILLER_35_780 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_22_441 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6878_ _7534_/Q _6878_/A2 _6879_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_50_761 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_139_148 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5829_ hold773/Z _5840_/A2 _5830_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_22_463 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_163_641 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_162_140 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_135_354 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_118_31 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_2_802 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_78_46 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_1_312 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
Xhold670 _7612_/Q hold670/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
Xhold681 hold681/I _7692_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
Xhold692 _7995_/I hold692/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
XFILLER_89_496 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_77_636 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_76_124 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_49_338 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_94_67 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_91_105 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_76_179 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_45_511 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_94_89 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_85_691 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_18_747 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_72_363 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_32_227 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_25_290 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_9_423 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_41_783 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_173_416 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_13_496 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_139_682 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_138_170 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_126_321 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xoutput208 _3703_/ZN mgmt_gpio_oeb[9] VDD VSS gf180mcu_fd_sc_mcu7t5v0__buf_4
Xoutput219 _7993_/Z mgmt_gpio_out[19] VDD VSS gf180mcu_fd_sc_mcu7t5v0__buf_4
XFILLER_175_70 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_154_685 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_107_590 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_4_183 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_141_357 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_68_614 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4160_ _7653_/Q _6022_/A1 hold194/I _7348_/Q _4779_/A1 _7477_/Q _4162_/A2 VDD VSS
+ gf180mcu_fd_sc_mcu7t5v0__aoi222_1
XFILLER_110_744 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4091_ _7638_/Q _5988_/A1 _4091_/B _4092_/A4 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_110_788 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_95_499 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_82_105 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7850_ hold61/Z _7877_/RN _7877_/CLK hold59/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_36_522 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6801_ _7107_/A1 _6767_/C _7433_/Q _6802_/B2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_63_352 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_63_341 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_24_717 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_7781_ _7781_/D _7877_/RN _7851_/CLK _7781_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
X_4993_ _5741_/A1 _5603_/A1 _4993_/B _4993_/C _4998_/C VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XFILLER_177_700 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_149_413 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6732_ _7923_/Q _7133_/S _6733_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_3944_ _7892_/Q _6520_/A1 _4488_/A1 _7361_/Q hold43/I _7746_/Q _3948_/A1 VDD VSS
+ gf180mcu_fd_sc_mcu7t5v0__aoi222_2
XFILLER_23_19 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_176_210 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_149_424 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3875_ _3886_/A2 hold82/Z _6384_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_4
X_6663_ _7910_/Q _7909_/Q _7908_/Q _6663_/A4 _6893_/C1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor4_4
XFILLER_177_777 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_176_265 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5614_ _5614_/A1 _5642_/A2 _5614_/A3 _5614_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__and3_1
XFILLER_31_282 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_176_276 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_136_118 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6594_ _6586_/B _6594_/A2 _7910_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_5545_ _5662_/A1 _5545_/A2 _5545_/B _5764_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi21_2
XFILLER_145_641 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_172_460 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5476_ _5527_/A1 _5498_/A2 _5476_/B _5523_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_145_696 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_117_354 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7215_ _4376_/B _7511_/Q _7941_/Q _7215_/C _7216_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai211_1
X_4427_ _7413_/Q _4427_/A2 _4427_/B _4428_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_132_368 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7146_ _7837_/Q _7203_/A2 _7193_/B1 _7635_/Q _7148_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_171_17 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_160_699 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_100_210 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_99_783 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_86_433 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4358_ _7432_/Q _7581_/Q _4359_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_58_124 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4289_ _7344_/Q _3734_/Z _7344_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_7077_ _7077_/A1 _7077_/A2 _7077_/A3 _7077_/A4 _7078_/A4 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand4_1
XFILLER_104_33 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_101_799 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6028_ _4460_/Z _6038_/A2 _6028_/B _7654_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_58_179 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_2105 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2116 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2149 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2138 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2127 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1415 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1404 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_70_812 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_64_59 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_64_37 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_27_566 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7979_ _7979_/D _7332_/Z _4415_/A2 _7979_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_2
XFILLER_120_21 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1448 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1437 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1426 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_81_171 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_14_205 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_54_396 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_120_65 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_120_54 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1459 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_168_744 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_10_400 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_23_761 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_23_783 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_168_788 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_109_800 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_148_490 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_108_321 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_89_34 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_136_663 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_97_709 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_123_357 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_2_676 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_150_176 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_145_73 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_77_499 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_64_105 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_18_522 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_73_672 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_45_352 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1960 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_158_210 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1993 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1982 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1971 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_9_231 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_174_747 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_3660_ _3660_/I _4370_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_9_286 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_139_490 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_127_641 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_161_419 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5330_ _5200_/B _3727_/I _5369_/B _5648_/B2 _5335_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand4_1
X_5261_ _5200_/B _3727_/I _5338_/A1 _5369_/B _5504_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand4_4
XFILLER_141_110 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_4212_ hold609/I _4212_/A2 _5849_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_48_2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7000_ _6949_/I _6997_/Z _7000_/A3 _7000_/A4 _7001_/B2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand4_1
X_5192_ _5200_/B _5230_/A1 _5663_/A1 _5371_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor3_1
XFILLER_141_165 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_141_176 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4143_ hold38/Z _3828_/I _4831_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_4074_ _3828_/I hold149/Z _5874_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_2
XFILLER_95_274 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_83_425 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_110_596 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_7902_ _7902_/D _7938_/RN _7940_/CLK _7902_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_55_138 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_70_108 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_52_812 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7833_ _7833_/D _7901_/RN _7833_/CLK _7833_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
X_7764_ _7764_/D _7877_/RN _7773_/CLK _7764_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
X_4976_ _4993_/B _5604_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_6715_ _7760_/Q _6892_/A2 _6893_/C1 _7630_/Q _6716_/A4 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_177_552 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_149_243 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_7695_ _7695_/D _7923_/RN _7735_/CLK _7695_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
X_3927_ _7940_/Q _7579_/Q _7580_/Q _3927_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_165_725 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3858_ hold89/Z hold54/Z _6282_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_4
X_6646_ _7910_/Q _6662_/A3 _6661_/A3 _6885_/B1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor3_4
XFILLER_50_17 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_3789_ _7337_/Q _7336_/Q _7414_/Q _3789_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_6577_ _7434_/Q _6590_/A1 _6586_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_5528_ _3727_/I _5528_/A2 _5552_/A4 _5540_/B2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor3_2
XFILLER_133_611 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_117_140 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_106_803 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_160_463 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5459_ _5752_/B1 _5668_/A2 _5459_/B _5668_/B _5460_/A4 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XFILLER_105_357 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_79_709 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_132_176 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_115_21 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_99_580 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_87_753 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_86_230 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7129_ _7129_/A1 _7129_/A2 _7129_/A3 _7128_/Z _7130_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand4_1
XFILLER_46_105 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_59_499 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_46_127 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_62_609 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1223 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1212 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1201 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_152_2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_91_35 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1256 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1245 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1234 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_168_530 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1289 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1278 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1267 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_399 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_168_585 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_156_747 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_171_706 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_109_641 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_10_274 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_6_256 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_170_238 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_123_110 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_163_290 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_151_430 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_69_208 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_151_496 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_97_528 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_77_241 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_49_70 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_93_712 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_65_447 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_65_425 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_93_767 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_92_266 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_1_99 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_34_812 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_52_108 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4830_ _7230_/A1 _4828_/S _4830_/B _7503_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
XTAP_1790 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_4761_ hold47/Z _4763_/A2 _4761_/B _7468_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_4692_ _3819_/Z _4454_/Z _4693_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_3712_ _7609_/Q _7107_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_6500_ _4481_/I _6502_/A2 _6500_/B _7876_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_7480_ _7480_/D _7949_/CLK _7480_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_3643_ hold52/Z _3801_/I0 VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_6431_ hold283/Z _6434_/A2 _6432_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_134_408 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6362_ _4476_/I _6366_/A2 _6362_/B hold236/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_155_780 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5313_ _5687_/C _5495_/B2 _5741_/B _5316_/C VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_142_463 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6293_ hold732/Z _6298_/A2 _6294_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_114_143 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_114_176 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_102_327 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5244_ _5779_/A1 _5433_/C _5273_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
Xhold18 hold18/I hold18/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
Xhold29 hold29/I hold29/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
X_5175_ _5749_/A2 _5175_/A2 _5178_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_96_561 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_28_105 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4126_ hold54/Z _3869_/I _4594_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_2
X_4057_ _4057_/A1 _4057_/A2 _4057_/A3 _4057_/A4 _4058_/A4 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand4_1
XFILLER_45_17 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_56_458 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_71_428 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_25_812 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_306 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
X_7816_ _7816_/D _7923_/RN _7816_/CLK _7816_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffsnq_1
XFILLER_101_34 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_339 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_328 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_317 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_51_141 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7747_ hold3/Z _7877_/RN _7747_/CLK _7747_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
X_4959_ _5797_/B _4965_/B _5774_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_4
XFILLER_61_27 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_7678_ _7678_/D _7923_/RN _7737_/CLK _7678_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffsnq_1
XFILLER_138_747 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_6629_ _6634_/A1 _7906_/Q _6659_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_165_566 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_153_728 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_118_460 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_180_525 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_3_215 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_180_558 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_145_290 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_161_783 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_133_496 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_133_485 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_105_176 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_160_282 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_121_658 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_120_179 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_86_57 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_75_712 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_59_252 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_59_274 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_19_73 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_47_425 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_142_63 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_142_52 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_47_458 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_16_812 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_27_160 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_34_108 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1031 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_130 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1020 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1064 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1053 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1042 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_129_703 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1097 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1086 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1075 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_185 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_30_347 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_11_561 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_51_82 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_137_780 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_124_463 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_804 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_815 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_826 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_97_347 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_837 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_848 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_859 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_85_509 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_25_4 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_93_531 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_65_211 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_65_200 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_65_266 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_53_406 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6980_ _7376_/Q _7188_/A2 _6990_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_5931_ hold340/Z _5936_/A2 hold341/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_25_119 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_53_428 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_80_247 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_34_620 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_179_647 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5862_ _4460_/Z _5868_/A2 _5862_/B hold388/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_33_141 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7601_ _7601_/D _7853_/RN _7601_/CLK _7601_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
X_5793_ _5104_/B _5793_/A2 _5793_/B _5794_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_4813_ hold409/Z _4816_/A2 hold410/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_178_179 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4744_ hold47/Z _4753_/S _4744_/B hold377/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_7532_ _7532_/D _7938_/RN _7532_/CLK _7532_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_147_522 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_119_224 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_119_246 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7463_ _7463_/D _7853_/RN _7600_/CLK _7463_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
X_4675_ _3879_/Z _4476_/I _4676_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_6414_ hold305/Z _6417_/A2 _6415_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_7394_ _7394_/D _7900_/RN _7767_/CLK _7394_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
X_6345_ _4476_/I _6349_/A2 _6345_/B hold344/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_1_708 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_143_783 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6276_ hold852/Z _6281_/A2 _6277_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
Xinput108 wb_adr_i[21] _5302_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__buf_3
X_5227_ _5199_/B _5201_/B _5338_/A1 _5369_/B _5573_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor4_4
XFILLER_130_433 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
Xinput119 wb_adr_i[31] _4367_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XFILLER_102_179 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_57_712 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5158_ _5496_/A1 _5527_/A1 _5167_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_84_531 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_29_425 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5089_ _3728_/I _5022_/B _5303_/A3 _5285_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand3_1
X_4109_ _4206_/A1 _7223_/A1 _4109_/B _4110_/I0 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_56_244 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_16_108 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_25_631 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_112_99 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_72_37 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_125 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_103 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_114 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_158 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_147 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_136 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_12_325 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_9_808 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_24_185 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_52_494 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_169 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_8_307 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_40_656 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_181_812 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_115_2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_106_463 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_121_444 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_94_306 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_153_73 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_121_499 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_47_200 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_63_704 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_48_756 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_35_428 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_90_534 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_62_247 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_47_299 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_15_141 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_5 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_30_188 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_172_812 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4460_ _4461_/A1 hold31/Z _4460_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__and2_4
XFILLER_156_385 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xhold307 _7788_/Q hold307/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
Xhold329 _7697_/Q hold329/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
Xhold318 hold318/I _7797_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
X_4391_ _4387_/S _7889_/Q _4391_/B _4391_/ZN VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_171_388 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_125_783 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_125_772 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_6130_ _4460_/Z _6140_/A2 _6130_/B hold643/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
XTAP_601 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_612 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_623 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_634 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_30_2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_97_144 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_6061_ hold652/Z _6072_/A2 _6062_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_645 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_656 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_667 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_58_509 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5012_ _4926_/Z _5010_/Z _5195_/B _5139_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_4
XTAP_678 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_689 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_39_712 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_66_542 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_66_531 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_38_266 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6963_ _7870_/Q _7195_/C1 _7207_/B1 _7716_/Q _6965_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_5914_ hold219/Z _5919_/A2 hold220/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_81_567 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6894_ _7400_/Q _6894_/A2 _6659_/Z _7471_/Q _6894_/C1 _7404_/Q _6895_/A4 VDD VSS
+ gf180mcu_fd_sc_mcu7t5v0__aoi222_1
X_5845_ _4454_/Z _5845_/A2 _5845_/B _7570_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_179_499 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_166_105 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_21_144 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_5776_ _5776_/A1 _5778_/A1 _5776_/A3 _5776_/A4 _5777_/C VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand4_1
X_7515_ _7515_/D _7959_/RN _7959_/CLK _7515_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_163_812 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_147_352 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_147_330 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_108_717 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_4727_ _6545_/A1 _4731_/A2 _4727_/B hold143/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_4658_ _7425_/Q _4685_/A1 _4661_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_7446_ _7446_/D _7900_/RN _7892_/CLK _8006_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
Xhold830 _7807_/Q hold830/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
XFILLER_135_558 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_123_709 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xinput90 spimemio_flash_io2_oeb input90/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyb_1
X_7377_ _7377_/D _7877_/RN _7381_/CLK _7377_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffsnq_1
Xhold852 _7771_/Q hold852/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
XFILLER_89_601 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
Xhold841 _7355_/Q hold841/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
Xhold863 _7374_/Q hold863/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
X_4589_ _4589_/A1 _6537_/A2 _4593_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_6328_ _4476_/I _6332_/A2 _6328_/B hold374/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_107_33 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xhold874 _7863_/Q hold874/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
Xhold885 _7613_/Q hold885/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
Xhold896 _7823_/Q hold896/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
XFILLER_131_775 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_131_764 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6259_ hold726/Z _6264_/A2 _6260_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_103_499 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_76_317 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_17_428 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_72_534 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_44_247 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_40_420 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_9_638 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_172_108 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_153_311 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_126_536 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_126_514 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_5_800 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_4_321 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_141_517 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_107_783 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_106_260 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_122_742 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_79_144 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_79_199 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_593 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_48_531 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_57_70 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_57_81 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_63_556 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_63_545 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_35_236 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_63_567 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3960_ hold609/Z _3959_/Z _4719_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_4
XFILLER_44_770 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3891_ _7619_/Q _5937_/A1 _4488_/A1 _7362_/Q _3892_/A4 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_5630_ _5776_/A1 _5778_/A1 _5697_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_31_486 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_148_149 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_5561_ _5741_/A1 _4993_/B _5663_/A1 _5561_/B _5562_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai31_1
XFILLER_78_2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7300_ _7901_/RN _4334_/Z _7300_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_145_812 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_144_311 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_5492_ _5648_/A1 _5735_/A2 _5685_/B _5648_/B2 _5642_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_4512_ hold285/Z _4521_/A2 hold286/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_7231_ _7281_/A2 _3658_/I _7233_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_172_664 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_117_558 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
Xhold115 hold115/I _7679_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
XFILLER_105_709 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xhold126 hold126/I _7703_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
Xhold104 _7769_/Q hold104/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
XFILLER_7_170 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_171_141 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4443_ hold21/I hold4/Z hold49/I hold5/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_4
Xhold148 _3803_/Z hold148/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
Xhold159 hold159/I _7821_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
XFILLER_132_528 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xhold137 _7619_/Q hold137/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
X_4374_ _4906_/S _4374_/A2 _4374_/A3 _4374_/A4 _4375_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand4_1
X_7162_ _7525_/Q _7190_/C1 _7168_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_6113_ _4460_/Z _6123_/A2 _6113_/B hold629/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_113_753 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7093_ _7891_/Q _7196_/A2 _7196_/B1 _7641_/Q _7095_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XTAP_442 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_431 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_420 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_6044_ hold678/Z _6055_/A2 _6045_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_140_594 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_464 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_475 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_453 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_100_458 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_497 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_486 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_82_810 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2309 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_7995_ _7995_/I _7995_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_54_534 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1619 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1608 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_6946_ _6946_/A1 _6946_/A2 _6946_/A3 _6946_/A4 _6946_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__and4_1
XFILLER_26_258 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_53_17 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6877_ _7133_/S _6877_/A2 _6877_/B _7929_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_167_436 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_167_425 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5828_ hold150/Z _6537_/A2 _5840_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_4
X_5759_ _5759_/A1 _5768_/A3 _5779_/A2 _5779_/A1 _5759_/C _5760_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi221_1
XFILLER_154_108 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_148_672 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_136_812 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7429_ _7429_/D _7923_/RN _7698_/CLK _7986_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_118_87 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_104_742 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
Xhold671 _7840_/Q hold671/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
XFILLER_78_25 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
Xhold660 _7642_/Q hold660/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
Xhold693 hold693/I _7421_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
Xhold682 _7800_/Q hold682/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
XFILLER_1_357 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_182_2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_134_97 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_18_737 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_27_73 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_27_95 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_33_718 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_45_567 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_60_548 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_13_442 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_13_453 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_40_250 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_158_458 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_173_428 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
Xclkbuf_3_7__f_csclk clkbuf_0_csclk/Z clkbuf_3_7__f_csclk/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_138_160 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_5_641 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_181_450 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_153_163 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_153_141 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_141_303 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xoutput209 _4405_/Z mgmt_gpio_out[0] VDD VSS gf180mcu_fd_sc_mcu7t5v0__buf_4
XFILLER_175_93 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_99_228 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_95_423 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_95_456 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4090_ _4090_/A1 _4090_/A2 _4090_/A3 _4091_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_36_534 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_48_383 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6800_ _6800_/A1 _6800_/A2 _6800_/A3 _6799_/Z _6802_/B1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand4_1
X_4992_ _5254_/A2 _5608_/A1 _4993_/C VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_4
X_7780_ _7780_/D _7853_/RN _7812_/CLK _7780_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_23_217 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_177_712 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6731_ _7433_/Q _7922_/Q _6731_/B1 _6731_/B2 _6733_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_3943_ _3943_/A1 _3943_/A2 _3943_/A3 _3943_/A4 _3954_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand4_2
X_6662_ _7910_/Q _6663_/A4 _6662_/A3 _6892_/B1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor3_4
X_3874_ hold42/Z hold82/Z _6333_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_4
X_5613_ _5359_/B _5613_/A2 _5678_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_136_108 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_118_812 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6593_ _7434_/Q _6767_/C _6593_/B1 _7910_/Q _6594_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_5544_ _5547_/A1 _5547_/A2 _5651_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_144_130 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5475_ _5066_/Z _5680_/A1 _5475_/B _5502_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_7214_ _7214_/A1 _7214_/A2 _7517_/D _7216_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_144_174 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4426_ _7412_/Q _7415_/Q _4427_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_7145_ _7829_/Q _7202_/A2 _7205_/B1 _7747_/Q _7148_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_98_250 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_101_712 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_101_701 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_100_200 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xclkbuf_leaf_93_csclk _7407_/CLK _7874_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
X_4357_ _7433_/Q _4361_/A2 _4359_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_4288_ _7345_/Q _4288_/A2 _7345_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__xnor2_1
X_7076_ _7818_/Q _7207_/A2 _7207_/B1 _7720_/Q _7076_/C _7077_/A4 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi221_1
XFILLER_104_12 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_101_778 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6027_ hold653/Z _6038_/A2 _6028_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_55_810 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2106 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2117 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2139 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2128 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1405 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_82_673 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7978_ _7978_/D _7331_/Z _4398_/I1 _7978_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XTAP_1438 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1427 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1416 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_81_150 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xclkbuf_leaf_31_csclk _7422_/CLK _7853_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_120_33 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1449 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_6929_ _6953_/A1 _6950_/A1 _6941_/A2 _7189_/C1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor3_4
XFILLER_168_734 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_120_99 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_80_37 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_22_250 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_155_428 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_109_812 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_182_247 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xclkbuf_leaf_46_csclk clkbuf_3_7__f_csclk/Z _7461_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_136_653 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_129_75 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_13_97 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_89_68 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_8_2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_2_600 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
Xhold490 _7628_/Q hold490/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
XFILLER_89_272 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_77_412 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_49_125 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_58_670 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_161_73 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_161_51 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_64_128 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_18_512 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_18_534 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_159_712 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1961 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1950 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_60_334 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_158_200 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1994 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1983 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1972 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_60_389 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_41_570 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_13_283 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_146_417 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_118_108 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_173_247 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_142_601 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5260_ _5199_/B _5201_/B _3728_/I _5022_/B _5768_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor4_4
XFILLER_141_144 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4211_ hold89/I _4075_/B _5855_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_5191_ _5476_/B _5689_/A2 _5191_/B1 _5191_/B2 _7520_/Q _5362_/B1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai221_1
XFILLER_110_531 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_110_520 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4142_ _7677_/Q _6073_/A1 _4174_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_68_478 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_4073_ _4427_/B _4073_/A2 _4073_/A3 _4073_/B hold941/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai31_1
XFILLER_110_586 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7901_ _7901_/D _7901_/RN _7901_/CLK _7901_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_95_286 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_55_128 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7832_ _7832_/D _7901_/RN _7901_/CLK _7832_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffsnq_1
XFILLER_64_673 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_169_509 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4975_ _5069_/A2 _4930_/Z _4953_/Z _4975_/A4 _4993_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand4_4
X_7763_ _7763_/D _7877_/RN _7773_/CLK _7763_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
X_6714_ _7816_/Q _6880_/A2 _6891_/B1 _7670_/Q _6716_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_3926_ hold149/Z _4155_/A2 _5870_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_4
XFILLER_51_389 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_7694_ _7694_/D _7853_/RN _7720_/CLK _7694_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffsnq_1
XFILLER_137_428 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6645_ _7910_/Q _6664_/A3 _6658_/A3 _6882_/B1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor3_4
X_3857_ _4075_/B _4217_/A2 hold194/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_4
XFILLER_164_247 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3788_ _3810_/S hold88/Z _3788_/B _3925_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi21_4
X_6576_ _6634_/A1 _6633_/A2 _6658_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_4
X_5527_ _5527_/A1 _5689_/A2 _5548_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_5458_ _5496_/A1 _5527_/A1 _5458_/B _5458_/C _5668_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi211_2
XFILLER_132_144 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_182_28 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_132_166 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_99_570 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5389_ _5705_/A2 _5585_/A1 _5624_/B _5759_/A1 _5736_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_4409_ input1/Z _7607_/Q _4409_/B _4409_/ZN VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_115_44 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_113_380 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_101_531 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7128_ _6949_/I _7128_/A2 _7128_/A3 _7128_/A4 _7128_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__and4_1
XFILLER_59_434 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_115_88 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_86_264 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_7059_ _7680_/Q _7191_/A2 _7190_/B1 _7616_/Q _7190_/A2 _7794_/Q _7063_/A1 VDD VSS
+ gf180mcu_fd_sc_mcu7t5v0__aoi222_1
XFILLER_74_459 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_43_802 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1213 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1202 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_27_364 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_1257 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1246 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1235 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1224 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_70_632 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_15_559 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_145_2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1279 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1268 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_70_676 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_42_356 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_42_389 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_23_570 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_168_575 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_128_417 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_155_247 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_11_798 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_124_601 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_108_141 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_170_228 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_170_217 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_124_667 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_123_144 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_151_486 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_2_463 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_77_231 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_77_286 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_19_810 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_92_245 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_92_234 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_18_342 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_92_278 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_65_81 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_65_70 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_46_673 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1780 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1791 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_4760_ hold587/Z _4763_/A2 _4761_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_146_203 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4691_ _7437_/Q _4718_/A1 _4694_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_119_428 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3711_ _7608_/Q _7079_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_81_91 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_174_534 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_146_247 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3642_ hold40/I _5640_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_6430_ _6549_/A1 _6434_/A2 _6430_/B _7843_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_6361_ hold235/Z _6366_/A2 _6362_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_60_2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5312_ _5724_/B _5624_/A2 _5741_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_6292_ _6547_/A1 _6298_/A2 _6292_/B _7778_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_114_155 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_102_317 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5243_ _5714_/B1 _5687_/B _5247_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_2
Xhold19 hold19/I hold19/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
XFILLER_130_648 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5174_ _5735_/A2 _5643_/A2 _5027_/Z _5643_/B1 _5175_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_69_732 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4125_ hold54/Z _3881_/Z _4554_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_56_404 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_110_394 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_84_735 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_83_212 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_69_798 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4056_ _7623_/Q _5954_/A1 _5988_/A1 _7639_/Q _4057_/A4 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XPHY_307 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_101_24 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_101_13 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_64_481 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7815_ _7815_/D _7923_/RN _7815_/CLK _7815_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffsnq_1
XPHY_329 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_318 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_52_676 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4958_ _4941_/C _4941_/B _4973_/A3 _4920_/Z _4965_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai22_4
X_7746_ _7746_/D _7877_/RN _7849_/CLK _7746_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_24_389 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_177_28 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_131_8 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3909_ _7354_/Q hold194/I _6124_/A1 _7707_/Q _3911_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_7677_ _7677_/D _7938_/RN _7738_/CLK _7677_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffsnq_1
X_4889_ hold768/Z _4892_/A2 _4890_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_138_759 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_137_225 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6628_ _7921_/Q _7133_/S _6686_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_117_6 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_4_717 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6559_ _7902_/Q _6559_/A2 _6560_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_145_280 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_106_667 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_106_656 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_105_144 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_160_250 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_120_103 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_79_529 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_120_158 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_120_147 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_86_69 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_59_264 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_59_286 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_47_415 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_28_673 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1010 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1021 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_70_440 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1065 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1054 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1032 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1043 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_35_73 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_1098 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1087 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1076 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_175 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_175_309 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_156_534 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_128_247 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_7_566 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_143_228 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_109_494 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_112_615 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_805 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_816 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_151_294 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_151_283 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_3_783 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_2_260 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_827 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_838 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_849 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_120_670 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_93_521 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5930_ _6547_/A1 _5936_/A2 _5930_/B hold541/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_7600_ hold20/Z _7923_/RN _7600_/CLK hold18/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_61_440 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5861_ _7577_/Q _5868_/A2 _5862_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_33_153 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_34_676 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5792_ hold52/I _5520_/C _5792_/B1 _5792_/B2 _5806_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_4812_ _4812_/A1 _7285_/A2 _4816_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_21_304 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4743_ hold375/Z _4753_/S hold376/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_7531_ _7531_/D _7938_/RN _7531_/CLK _7531_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
X_7462_ _7462_/D _7853_/RN _7600_/CLK _7462_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
X_4674_ hold612/Z _4685_/A1 _4677_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_6413_ _6549_/A1 _6417_/A2 _6413_/B _7835_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_134_206 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_128_770 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7393_ _7393_/D _7900_/RN _7881_/CLK _7393_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
X_6344_ hold343/Z _6349_/A2 _6345_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_163_19 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_142_250 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6275_ _6547_/A1 _6281_/A2 _6275_/B _7770_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
Xinput109 wb_adr_i[22] _5224_/A4 VDD VSS gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_170_592 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5226_ _5006_/C _5616_/A1 _5433_/C _5290_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_130_489 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5157_ _5179_/B _5783_/A2 _5173_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_5088_ _5338_/A1 _5369_/B _5054_/Z _5114_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor3_2
XFILLER_96_392 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4108_ _7549_/Q _4206_/A1 _4109_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_56_256 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_57_768 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_71_215 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_4039_ _4039_/I0 hold949/Z _4427_/B _7552_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_112_45 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_25_621 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_72_49 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_40_602 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_104 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_115 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_148 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_137 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_126 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
X_7729_ _7729_/D _7877_/RN _7729_/CLK _7729_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XPHY_159 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_138_534 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_20_392 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_125_228 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_108_2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_180_389 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_161_570 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_140_209 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_137_97 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_133_283 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_764 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_87_392 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_47_223 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XPHY_6 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_16_676 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_16_665 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_62_60 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_156_342 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_129_567 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_144_526 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_144_515 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
Xhold308 hold308/I _7788_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
XFILLER_7_77 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4390_ _4387_/S input90/Z _4391_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
Xhold319 _7354_/Q hold319/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
XFILLER_171_367 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_124_250 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_98_624 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_98_602 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_98_635 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_602 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_613 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_624 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_635 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_646 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_657 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_668 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_6060_ _4454_/Z _6072_/A2 _6060_/B _7669_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_5011_ _5211_/A3 _5011_/A2 _5011_/B _5016_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi21_2
XFILLER_78_370 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_23_2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_679 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_78_392 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_38_245 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_66_587 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6962_ _7894_/Q _7197_/A2 _7189_/C1 _7652_/Q _6965_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_53_215 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_53_237 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5913_ hold16/Z _5919_/A2 hold19/Z hold20/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_22_602 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6893_ _7402_/Q _6893_/A2 _6893_/B1 _7390_/Q _6893_/C1 _7473_/Q _6895_/A3 VDD VSS
+ gf180mcu_fd_sc_mcu7t5v0__aoi222_1
X_5844_ hold897/Z _5845_/A2 _5845_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_22_646 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_166_139 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7514_ _7514_/D _7959_/RN _7545_/CLK _7514_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
X_5775_ _5775_/A1 _5775_/A2 _5801_/A1 _5786_/C1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand3_1
X_4726_ hold141/Z _4731_/A2 hold142/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_4657_ _4685_/A1 _4657_/A2 _4657_/B hold516/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_7445_ _7445_/D _7875_/RN _7881_/CLK _7445_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
X_7376_ _7376_/D _7877_/RN _7381_/CLK _7376_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffsnq_1
XFILLER_162_334 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
Xinput91 spimemio_flash_io3_do input91/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyb_1
Xinput80 spi_sck input80/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyb_1
Xhold820 hold820/I _4882_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
Xhold831 _7749_/Q hold831/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
XFILLER_162_389 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xhold864 _7375_/Q hold864/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
X_6327_ hold372/Z _6332_/A2 hold373/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
Xhold842 hold842/I _4490_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
Xhold853 _7467_/Q hold853/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
X_4588_ _4454_/Z _4588_/A2 _4588_/B _7398_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_143_570 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_115_294 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_115_283 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_107_45 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_88_123 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
Xhold875 _7799_/Q hold875/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
Xhold897 _7570_/Q hold897/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
Xhold886 _7524_/Q hold886/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
XFILLER_131_754 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6258_ _6547_/A1 _6264_/A2 _6258_/B _7762_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_77_808 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5209_ _5209_/A1 _5209_/A2 _5209_/A3 _5376_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand3_2
X_6189_ hold233/Z _6191_/A2 _6189_/B _7730_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_131_798 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_97_690 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_29_212 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_69_392 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_29_245 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_57_543 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_57_554 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_13_635 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_12_134 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_8_105 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_166_673 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_5_812 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_32_96 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_181_665 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_106_250 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_180_186 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_121_231 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_121_286 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_121_275 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_95_638 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_94_126 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_79_189 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_94_159 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_35_204 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_90_321 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_35_215 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_73_70 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_149_618 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_3890_ _7382_/Q hold55/I _6452_/A1 _7861_/Q _3892_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_31_432 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5560_ _5613_/A2 _5560_/A2 _5590_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_5491_ _5542_/A2 _5542_/A3 _5517_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_8_672 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4511_ _4460_/Z _4521_/A2 _4511_/B hold633/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_4442_ hold21/Z _3810_/S _4442_/B hold22/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi21_4
Xhold116 _7671_/Q hold116/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
Xhold105 hold105/I _7769_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
X_7230_ _7230_/A1 _7228_/S _7230_/B _7949_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_7_160 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_172_676 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_171_164 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
Xhold138 hold138/I _7619_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
Xhold127 _7655_/Q hold127/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
XFILLER_104_209 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xhold149 hold149/I hold149/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
X_4373_ _4925_/A1 _4923_/A1 _4365_/Z _4374_/A4 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor3_1
XFILLER_144_389 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_125_570 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7161_ _7133_/S _7161_/A2 _7161_/A3 _7161_/B _7938_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai31_1
X_6112_ hold627/Z _6123_/A2 hold628/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_113_776 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_86_605 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7092_ _7649_/Q _7195_/A2 _7195_/B1 _7625_/Q _7195_/C1 _7875_/Q _7097_/A3 VDD VSS
+ gf180mcu_fd_sc_mcu7t5v0__aoi222_1
XFILLER_59_808 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_432 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_421 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_410 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_6043_ _4454_/Z _6055_/A2 _6043_/B _7661_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_85_104 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_465 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_476 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_454 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_443 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_58_318 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_85_148 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_498 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_487 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_7994_ _7994_/I _7994_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_1609 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_81_354 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6945_ _7189_/C1 _7190_/B1 _7196_/A2 _7193_/C1 _6946_/A4 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor4_1
XFILLER_35_760 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_179_231 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_81_398 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_35_771 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_41_207 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6876_ _7929_/Q _7133_/S _6877_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_179_286 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_10_605 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5827_ _6547_/A1 _5827_/A2 _5827_/B _7562_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_5758_ _5614_/Z _5758_/A2 _5758_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_182_418 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4709_ hold219/Z _3819_/Z _4709_/B _4710_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_135_312 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5689_ _5689_/A1 _5689_/A2 _5757_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_7428_ _7428_/D _7923_/RN _7597_/CLK _7985_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
Xhold661 _7714_/Q hold661/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
XFILLER_78_37 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xhold650 hold650/I _4515_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
Xhold672 _7732_/Q hold672/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
X_7359_ _7359_/D input75/Z _7570_/CLK _7359_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
Xhold694 _7776_/Q hold694/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
Xhold683 _7832_/Q hold683/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
XFILLER_89_443 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_134_32 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_103_275 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_77_638 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_134_54 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_103_286 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_175_2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_72_321 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_17_215 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_57_384 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_33_708 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_60_538 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_26_782 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_9_425 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_43_73 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_159_73 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_158_448 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_145_109 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_154_676 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_153_175 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_107_570 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_4_34 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_68_605 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_4_45 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_122_595 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_91_641 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_90_140 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_63_354 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4991_ _5206_/A2 _5136_/A1 _5585_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_4
X_6730_ _7027_/A1 _6767_/C _7433_/Q _6731_/B2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_90_195 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3942_ _7353_/Q hold194/I _4249_/A2 input32/Z _3943_/A4 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_176_212 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3873_ hold72/Z _4141_/A1 _6107_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_4
XFILLER_90_2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_32_763 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_32_774 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6661_ _6878_/A2 _6662_/A3 _6661_/A3 _6894_/C1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor3_4
X_5612_ _5599_/Z _5612_/A2 _5610_/Z _5639_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand3_1
X_6592_ _6618_/A3 _6830_/B _6593_/B1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_164_407 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5543_ _5741_/A3 _5545_/A2 _5543_/B _5543_/C _5547_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XFILLER_117_312 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_144_142 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_5474_ _5461_/Z _5474_/A2 _5474_/B _5521_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_117_378 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_132_326 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7213_ _7133_/S _7213_/A2 _7213_/B _7940_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_4425_ _7979_/Q _4425_/A2 _4425_/ZN VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_7144_ _7140_/Z _7144_/A2 _7144_/A3 _7144_/A4 _7159_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand4_1
XFILLER_99_763 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_4356_ _6937_/A1 _6953_/A1 _6950_/A1 _4361_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor3_1
XFILLER_59_638 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4287_ _7346_/Q _4287_/A2 _7346_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XFILLER_140_392 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_101_757 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_100_212 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7075_ _7075_/A1 _7075_/A2 _7075_/A3 _7076_/C VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_101_768 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6026_ _4454_/Z _6038_/A2 _6026_/B _7653_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
XTAP_2107 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_67_693 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_67_682 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_54_321 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2129 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2118 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1406 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_15_708 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7977_ _7977_/D _7330_/Z _4415_/A2 _7977_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XTAP_1439 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1428 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1417 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_538 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6928_ _7914_/Q _7913_/Q _6937_/A1 _6599_/Z _7200_/B1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor4_4
XFILLER_167_212 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_80_27 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_10_402 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_23_763 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6859_ _6859_/A1 _6859_/A2 _6859_/A3 _6860_/C VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_50_560 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_6_417 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_136_676 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_108_389 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_151_657 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_150_156 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xhold480 hold480/I _5851_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
Xhold491 _7598_/Q hold491/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
XFILLER_1_144 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_49_148 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_77_479 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_58_660 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_45_321 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_58_682 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_73_641 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_45_354 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_73_674 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_33_527 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_33_516 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_33_505 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1951 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1940 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_158_212 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1995 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1984 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1973 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1962 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_60_379 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_173_215 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_158_278 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_173_226 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_173_237 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_167_790 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_126_142 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_141_101 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_127_698 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_5_472 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_142_668 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_142_646 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4210_ _7586_/Q _5881_/A1 _4754_/A1 _7466_/Q _4243_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_5190_ _5424_/A1 _5680_/B2 _5755_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_122_392 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_96_744 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4141_ _4141_/A1 _3959_/Z _4873_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_96_788 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_37_800 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4072_ hold940/Z _4427_/B _4073_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_7900_ _7900_/D _7900_/RN _7900_/CLK _7900_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_37_811 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_48_170 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_64_630 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_36_321 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_48_181 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_91_460 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_63_140 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_24_527 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_36_387 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7831_ _7831_/D _7875_/RN _7862_/CLK _7831_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffsnq_1
XFILLER_51_302 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4974_ _5201_/B _5210_/A3 _4974_/A3 _5797_/C VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand3_4
X_7762_ _7762_/D _7877_/RN _7869_/CLK _7762_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_24_538 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_149_212 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3925_ hold26/Z _3925_/A2 hold75/Z hold71/Z _4155_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand4_4
X_6713_ _7702_/Q _6889_/A2 _6887_/B1 _7678_/Q _6659_/Z _7622_/Q _6716_/A2 VDD VSS
+ gf180mcu_fd_sc_mcu7t5v0__aoi222_1
X_7693_ _7693_/D _7938_/RN _7733_/CLK _7693_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffsnq_1
XFILLER_51_357 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6644_ _7910_/Q _6665_/A2 _6659_/A3 _6644_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__and3_2
XFILLER_165_716 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3856_ _3783_/Z hold41/Z hold75/Z hold71/Z _4217_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand4_4
XFILLER_20_744 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3787_ hold40/Z hold88/I _3810_/S hold41/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_4
X_6575_ _7907_/Q _7906_/Q _6590_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_2
X_5526_ _5066_/Z _5680_/B2 _5552_/A4 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_118_676 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5457_ _5741_/A3 _5099_/B _5776_/A1 _3723_/I _5457_/C _5459_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai221_1
XFILLER_133_635 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4408_ input1/Z input2/Z _4409_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_120_318 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_99_582 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5388_ _5772_/A1 _5614_/A1 _5783_/C VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_59_413 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4339_ _7518_/Q _4438_/A2 _7513_/Q _4340_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_115_23 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7127_ _7754_/Q _7201_/A2 _7205_/B1 _7746_/Q _7128_/A4 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_115_56 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_7058_ _7133_/S _7058_/A2 _7058_/A3 _7058_/B _7934_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai31_1
XFILLER_86_254 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6009_ _4454_/Z _6021_/A2 _6009_/B _7645_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_55_641 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_82_460 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1214 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1203 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1247 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1236 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1225 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_54_195 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_1269 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1258 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_24_31 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_24_53 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_138_2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_155_215 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_6_258 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_6_247 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_156_52 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_112_808 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_104_392 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_78_744 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_93_703 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_78_788 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_1_13 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_49_83 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_18_321 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_73_460 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_179_808 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_60_110 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_178_318 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1770 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_33_357 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1781 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1792 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_81_70 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_60_176 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xclkbuf_leaf_92_csclk _7407_/CLK _7822_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
X_3710_ _7623_/Q _3710_/ZN VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_4690_ _4718_/A1 _4690_/A2 _4690_/B hold562/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_3641_ hold74/I _5522_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_146_259 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6360_ _6547_/A1 _6366_/A2 _6360_/B _7810_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_142_410 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5311_ _5645_/A1 _5687_/B _5624_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_4
XFILLER_53_2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_182_590 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_127_495 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6291_ hold589/Z _6298_/A2 _6292_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_114_123 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_130_605 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_102_307 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5242_ _5689_/A1 _5563_/B2 _5575_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_5173_ _5476_/B _5498_/A2 _5173_/B _5173_/C _5178_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_68_243 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4124_ _3828_/I hold82/Z _4579_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_110_362 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_84_747 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_68_298 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
Xinput1 debug_mode input1/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
Xclkbuf_leaf_45_csclk clkbuf_3_7__f_csclk/Z _7456_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
X_4055_ input38/Z _5903_/A1 _5971_/A1 _7631_/Q _4057_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_37_641 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_91_290 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_36_195 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_7814_ _7814_/D _7938_/RN _7815_/CLK _7814_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffsnq_1
XFILLER_169_318 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_319 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_308 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_101_36 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_24_368 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4957_ _5069_/A2 _4930_/Z _4953_/Z _4957_/A4 _5797_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand4_4
XFILLER_101_69 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7745_ _7745_/D _7853_/RN _7818_/CLK _7745_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_177_362 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3908_ _7747_/Q hold43/I _4232_/A2 input10/Z _3911_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_7676_ _7676_/D _7938_/RN _7738_/CLK _7676_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffsnq_1
X_4888_ _4888_/A1 _6537_/A2 _4892_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_137_215 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3839_ hold27/Z hold54/Z _6299_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_4
X_6627_ _6556_/B _7002_/B _7133_/S VDD VSS gf180mcu_fd_sc_mcu7t5v0__and2_4
X_6558_ _7433_/Q _4331_/Z _6562_/A1 _4352_/B _6564_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_2
XFILLER_106_602 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_10_11 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_5509_ _5509_/A1 _5509_/A2 _5505_/Z _5509_/A4 _5519_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor4_1
X_6489_ hold903/Z _6502_/A2 _6490_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_121_627 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_121_638 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_86_37 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_142_87 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_90_717 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_83_780 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_55_460 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_42_110 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_55_493 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1000 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1011 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1022 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_70_463 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_1055 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1033 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1044 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_15_346 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_15_357 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_31_806 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1099 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1088 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1077 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1066 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_187 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_128_204 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_167_73 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_51_73 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_152_730 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_112_605 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_97_305 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_3_773 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_2_250 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_806 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_817 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_828 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_839 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_111_137 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_93_511 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_78_585 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_66_747 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_65_224 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_19_641 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_46_460 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5860_ hold64/Z _5868_/A2 _5860_/B hold65/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_179_638 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4811_ _7230_/A1 _4809_/S _4811_/B _7493_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
XTAP_2290 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_5791_ _5691_/Z _5791_/A2 _5760_/Z _5791_/A4 _5792_/B2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand4_1
XFILLER_61_496 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_61_485 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_175_800 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_4742_ _3879_/Z _4742_/A2 _4753_/S VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_4
X_7530_ _7530_/D _7961_/RN _7961_/CLK _7530_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_174_321 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7461_ _7461_/D _7853_/RN _7461_/CLK _7461_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
X_4673_ _4685_/A1 _4673_/A2 _4673_/B hold383/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_119_215 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_135_708 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_119_248 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6412_ hold727/Z _6417_/A2 _6413_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_7392_ _7392_/D _7900_/RN _7823_/CLK _7392_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_89_806 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6343_ _6547_/A1 _6349_/A2 _6343_/B _7802_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_6274_ hold437/Z _6281_/A2 _6275_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_209 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_103_638 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_102_104 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5225_ _5563_/B2 _5687_/B _5624_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_4
XFILLER_130_457 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5156_ _5600_/A1 _5797_/B _5797_/A2 _5542_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor3_1
XFILLER_69_574 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5087_ _4898_/Z _5777_/A1 _5087_/B _5087_/C _5094_/B1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai211_1
X_4107_ _4107_/A1 _4107_/A2 _4107_/A3 _7223_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor3_4
XFILLER_37_460 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4038_ _4284_/A1 _4826_/A1 _4038_/B _4039_/I0 VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_65_780 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_25_611 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_13_806 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_105 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_116 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_149 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_138 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_127 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
X_5989_ hold825/Z _6004_/A2 _5990_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_12_327 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_24_176 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_52_463 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_178_671 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7728_ hold29/Z _7877_/RN _7729_/CLK _7728_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_40_669 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_165_354 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7659_ _7659_/D _7923_/RN _7735_/CLK _7659_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_180_335 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_137_87 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_97_69 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
Xoutput190 _3685_/ZN mgmt_gpio_oeb[27] VDD VSS gf180mcu_fd_sc_mcu7t5v0__buf_4
XFILLER_0_754 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_153_64 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_48_747 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_28_460 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_7 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_55_290 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_71_783 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_70_271 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_31_636 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_43_496 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_30_124 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_156_321 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_8_810 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_30_179 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_116_207 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xhold309 _7877_/Q hold309/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
XFILLER_109_281 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_171_357 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_140_733 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_112_413 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_3_570 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_603 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_614 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_625 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_5010_ _5200_/B _5201_/B _5230_/A1 _5024_/A2 _5010_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__or4_4
XTAP_636 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_647 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_658 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_669 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_16_2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_38_268 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_47_780 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6961_ _7822_/Q _7202_/A2 _7196_/B1 _7636_/Q _7196_/A2 _7886_/Q _6967_/A2 VDD VSS
+ gf180mcu_fd_sc_mcu7t5v0__aoi222_1
X_5912_ hold18/Z _5919_/A2 hold19/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_6892_ _7386_/Q _6892_/A2 _6892_/B1 _7532_/Q _6895_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_5843_ _6539_/A1 _5845_/A2 _5843_/B _7569_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_34_463 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_167_619 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_61_282 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7513_ _7513_/D _7959_/RN _7545_/CLK _7513_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
X_5774_ _5774_/A1 _5774_/A2 _5774_/B1 _5774_/B2 _5774_/C _5801_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi221_2
XFILLER_175_641 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_147_354 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_147_332 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4725_ _4460_/Z _4731_/A2 _4725_/B hold417/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_30_680 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_174_140 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_162_313 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4656_ hold375/Z _3879_/Z _4656_/B _4657_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_107_207 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_7444_ _7444_/D _7875_/RN _7881_/CLK _7444_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_174_195 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_174_19 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7375_ _7375_/D _7877_/RN _7381_/CLK _7375_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffsnq_1
Xinput70 mgmt_gpio_in[7] input70/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyc_1
Xinput81 spi_sdo input81/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyb_1
Xhold810 hold810/I _4857_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
Xhold821 hold821/I _7532_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
X_4587_ hold855/Z _4588_/A2 _4588_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_131_700 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6326_ _6547_/A1 _6332_/A2 _6326_/B _7794_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_116_763 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xinput92 spimemio_flash_io3_oeb input92/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XFILLER_89_603 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xhold843 hold843/I _7355_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
XFILLER_1_507 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
Xhold832 _7388_/Q hold832/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
Xhold854 _7822_/Q hold854/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
Xhold865 _7456_/Q hold865/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
Xhold898 _7356_/Q hold898/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
Xhold887 hold887/I _4862_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
Xhold876 _7879_/Q hold876/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
XFILLER_131_766 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6257_ hold588/Z _6264_/A2 _6258_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_67_28 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_67_17 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5208_ _5015_/B _5197_/Z _5392_/A2 _5709_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor3_2
X_6188_ hold397/Z _6191_/A2 _6189_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_88_179 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5139_ _5139_/A1 _5014_/Z _5209_/A1 _5498_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand3_2
XFILLER_84_396 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_25_463 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_53_783 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_12_124 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_25_496 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_9_629 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_138_321 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_12_179 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_32_53 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_153_313 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_120_2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_153_357 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_141_519 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_180_176 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_134_582 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_4_389 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_4_378 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_122_744 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_122_788 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_562 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_102_490 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_63_503 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_48_566 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_63_514 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_29_780 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_35_238 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_51_709 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_16_463 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_148_129 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_157_641 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_31_499 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5490_ _5543_/B _5498_/A2 _5497_/A3 _5542_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor3_1
XFILLER_129_354 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4510_ hold631/Z _4521_/A2 hold632/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_171_121 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4441_ hold4/Z hold49/I _4442_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__and2_1
Xhold106 _7573_/Q hold106/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
Xhold117 hold117/I _6064_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
X_7160_ _7611_/Q _7210_/A2 _7160_/B _7433_/Q _7161_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi211_1
Xhold128 _7735_/Q hold128/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
Xhold139 _7627_/Q hold139/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
X_4372_ _4372_/A1 _4372_/A2 _4372_/A3 _4372_/A4 _4375_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand4_1
XFILLER_171_176 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_98_411 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_400 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_6111_ _4454_/Z _6123_/A2 _6111_/B hold924/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_140_530 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7091_ _7697_/Q _7194_/A2 _7194_/B1 _7665_/Q _7194_/C1 _7811_/Q _7097_/A2 VDD VSS
+ gf180mcu_fd_sc_mcu7t5v0__aoi222_1
XTAP_433 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_422 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_411 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_6042_ hold890/Z _6055_/A2 _6043_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_140_585 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_113_799 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_455 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_466 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_444 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_100_449 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_100_438 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_499 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_488 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_477 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_39_522 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_82_812 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7993_ _7993_/I _7993_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_81_333 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6944_ _7195_/B1 _7194_/B1 _7203_/B1 _7200_/B1 _6946_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor4_1
XFILLER_22_400 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_35_783 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6875_ _7433_/Q _7928_/Q _6875_/B1 _6875_/B2 _6877_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_5826_ hold548/Z _5827_/A2 _5827_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_5757_ _5425_/B _5757_/A2 _5757_/B _5783_/B _5758_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi211_1
X_4708_ _3819_/Z _4476_/I _4709_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_135_302 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_163_633 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5688_ _5705_/B _5555_/B _5688_/A3 _5725_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor3_1
X_7427_ _7427_/D _7853_/RN _7603_/CLK _7984_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_163_666 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4639_ hold420/Z _3830_/Z _4639_/B _4640_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_135_357 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_118_45 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_162_176 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xhold662 hold662/I _6155_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
XFILLER_118_89 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_116_560 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
Xhold640 hold640/I _7734_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
Xhold651 hold651/I _7367_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
X_7358_ _7358_/D _7961_/RN _7570_/CLK _7358_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffsnq_1
Xhold684 _7848_/Q hold684/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
Xhold695 _7742_/Q hold695/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
XFILLER_104_755 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_104_744 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6309_ _6547_/A1 _6315_/A2 _6309_/B _7786_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_7289_ _4454_/Z _7289_/A2 _7289_/B _7961_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
Xhold673 hold673/I _6194_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
XFILLER_131_574 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_131_563 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_104_799 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_89_499 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_76_105 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_134_88 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_94_37 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_94_48 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_168_2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_150_32 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_84_193 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_9_415 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_41_764 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_139_641 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_13_499 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_43_85 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_173_408 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_159_85 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_154_666 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_181_496 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_175_73 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_141_349 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_122_585 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_110_747 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_95_425 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_82_108 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_64_812 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_75_171 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4990_ _5394_/A1 _5254_/A2 _5136_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_2
XFILLER_17_783 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_23_208 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3941_ _7852_/Q _6435_/A1 _6265_/A1 _7772_/Q _3943_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_3872_ _3886_/A2 _4141_/A1 _6124_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_4
X_6660_ _7910_/Q _6664_/A2 _6664_/A3 _6884_/B1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor3_4
XFILLER_177_769 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_5611_ _5672_/A2 _5606_/B _5749_/A4 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_83_2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6591_ _7910_/Q _6879_/A1 _6767_/C VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_4
X_5542_ _5166_/B _5542_/A2 _5542_/A3 _5542_/A4 _5542_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__or4_1
XFILLER_145_611 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_144_121 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_172_463 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_117_368 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_117_357 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5473_ _5473_/A1 _5473_/A2 _5776_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_144_176 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4424_ _4424_/A1 input73/Z _4424_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__and2_1
X_7212_ _7940_/Q _7133_/S _7213_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_7143_ _7813_/Q _7194_/C1 _7204_/A2 _7845_/Q _7144_/A4 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_4355_ _7912_/Q _6599_/A2 _6950_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_4
XFILLER_98_274 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_7074_ hold57/I _7201_/A2 _7201_/B1 _7672_/Q _7075_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_58_105 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4286_ _7345_/Q _7344_/Q _3734_/Z _4287_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_113_596 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_104_14 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6025_ hold926/Z _6038_/A2 _6026_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_2108 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_55_812 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2119 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_7976_ _7976_/D _7329_/Z _4398_/I1 _7976_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XTAP_1429 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1418 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1407 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_81_163 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_81_141 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6927_ _6950_/A1 _6955_/A4 _6908_/Z _7194_/C1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor3_4
XFILLER_120_79 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_23_775 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_23_753 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_6858_ _7494_/Q _6882_/B1 _6647_/Z _7468_/Q _6859_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_168_747 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5809_ _6539_/A1 _5811_/A2 _5809_/B _7546_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_148_460 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6789_ _7665_/Q _6885_/A2 _6647_/Z _7617_/Q _6887_/B1 _7681_/Q _6791_/A2 VDD VSS
+ gf180mcu_fd_sc_mcu7t5v0__aoi222_1
XFILLER_182_238 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_135_121 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_124_806 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_163_496 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_135_176 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_2_602 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_145_43 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_89_230 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
Xhold470 _7361_/Q hold470/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
Xhold481 hold481/I _7572_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
XFILLER_2_646 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_150_179 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_150_168 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_145_65 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xhold492 hold492/I _5909_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
XFILLER_145_98 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_77_425 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_77_469 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_64_108 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_46_812 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_18_536 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_159_703 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1952 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1941 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1930 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_72_196 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_26_580 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_26_591 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1985 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1974 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1963 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_41_561 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1996 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_9_212 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_174_717 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_158_268 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_127_633 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_115_806 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_182_772 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_154_463 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_126_176 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_126_198 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_79_70 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4140_ _3828_/I hold54/Z _4584_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_2
XFILLER_68_447 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_68_458 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4071_ _7550_/Q _4206_/A1 _4073_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_83_428 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7830_ _7830_/D _7875_/RN _7830_/CLK _7830_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffsnq_1
XFILLER_63_152 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4973_ _3727_/I _4920_/Z _4973_/A3 _4975_/A4 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor3_2
X_7761_ _7761_/D _7901_/RN _7833_/CLK _7761_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_36_399 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6712_ _7734_/Q _6878_/A2 _6712_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__or2_1
X_3924_ input9/Z _4232_/A2 _3940_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_7692_ _7692_/D _7938_/RN _7733_/CLK _7692_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffsnq_1
XFILLER_51_369 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_20_734 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6643_ _7910_/Q _6663_/A4 _6664_/A2 _6881_/B1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor3_4
X_3855_ hold27/Z hold82/Z _6435_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_4
X_3786_ hold49/Z hold40/Z _3788_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__and2_1
X_6574_ _6633_/A2 _6618_/A3 _6574_/B _7906_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_5525_ _5543_/C _5498_/B _5545_/A2 _5542_/A4 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor3_1
XFILLER_173_783 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5456_ _5087_/B _5456_/A2 _5433_/C _5457_/C VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_117_176 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_105_305 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_145_496 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_105_349 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4407_ _7607_/Q _4334_/Z _4407_/B _4407_/ZN VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_132_179 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_132_168 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5387_ _5600_/A1 _5797_/B _4993_/C _5618_/A3 _5409_/B2 _5587_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai32_1
XFILLER_87_712 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4338_ _5903_/A2 _4338_/A2 _4338_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__or2_1
X_7126_ _7820_/Q _7207_/A2 _7207_/B1 _7722_/Q _7205_/A2 _7738_/Q _7128_/A3 VDD VSS
+ gf180mcu_fd_sc_mcu7t5v0__aoi222_1
XFILLER_59_425 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7057_ _7934_/Q _7133_/S _7058_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_28_801 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4269_ _7862_/Q _6469_/A1 _6537_/A1 _7894_/Q _4271_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_6008_ hold882/Z _6021_/A2 _6009_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_46_108 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1204 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_70_601 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7959_ _7959_/D _7959_/RN _7959_/CLK hold4/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XTAP_1248 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1237 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1226 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1215 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_168_511 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1259 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_168_522 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_11_712 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_155_238 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_149_780 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_10_266 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_136_474 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_136_463 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_156_64 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_151_444 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_123_157 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_123_146 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_2_454 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_172_41 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_151_499 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_49_73 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_65_428 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_19_812 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_105_90 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_92_247 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_45_141 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_73_494 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1760 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1782 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1793 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1771 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_159_566 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_174_514 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_147_739 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3640_ hold70/I _5362_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_60_4 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_155_783 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_154_271 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_127_485 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6290_ _6545_/A1 _6298_/A2 _6290_/B _7777_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_5310_ _5687_/C _5495_/B2 _5550_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_170_731 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_154_282 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_142_422 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_103_809 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5241_ _5199_/B _5201_/B _4915_/Z _5422_/B _5623_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand4_2
XFILLER_114_168 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_69_712 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_46_2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5172_ _5669_/A1 _5027_/Z _5173_/C VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_114_179 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_96_531 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_122_190 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4123_ hold54/Z _4151_/A2 _4564_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_4054_ _7671_/Q _6056_/A1 hold43/I hold68/I _4057_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_84_726 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
Xinput2 debug_oeb input2/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XFILLER_28_108 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_37_620 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
Xclkbuf_opt_1_0_csclk clkbuf_3_3__f_csclk/Z clkbuf_opt_1_0_csclk/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_36_141 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7813_ _7813_/D _7853_/RN _7853_/CLK _7813_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XPHY_309 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
X_7744_ hold44/Z _7901_/RN _7849_/CLK _7744_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_24_358 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_51_144 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4956_ _4944_/Z _4956_/A2 _5602_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_2
XFILLER_51_166 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_138_717 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7675_ _7675_/D _7853_/RN _7818_/CLK _7675_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
X_3907_ input28/Z _4239_/A2 _6367_/A1 _7821_/Q _3911_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_4887_ _4454_/Z _4887_/A2 _4887_/B hold793/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_20_531 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3838_ hold53/Z _3864_/A2 _3843_/A3 _3864_/A4 hold54/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand4_4
X_6626_ _7001_/C _7434_/Q _7002_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_153_709 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_20_597 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6557_ _6557_/I _6559_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_3769_ hold62/I hold962/Z _3772_/S _7969_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_118_463 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5508_ _5765_/A2 _5508_/A2 _5649_/A3 _5509_/A4 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_145_271 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6488_ _6539_/A1 _6502_/A2 _6488_/B _7870_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_160_252 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_126_34 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5439_ _5727_/A2 _5439_/A2 _5439_/A3 _5439_/A4 _5445_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand4_1
XFILLER_160_274 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_133_499 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_126_56 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_120_105 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_87_531 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_120_149 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7109_ _7133_/S _7109_/A2 _7109_/B _7936_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_47_428 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_142_44 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_74_247 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_90_729 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_27_141 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1001 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1012 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_150_2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1056 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1034 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1045 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1023 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_70_486 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_70_475 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1089 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1078 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1067 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_35_97 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_30_339 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_156_514 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_137_783 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_109_463 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_152_742 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_136_271 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_109_496 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_152_753 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_807 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_818 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_829 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_78_531 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_93_567 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_93_589 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_34_601 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_61_420 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_178_105 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2280 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_33_144 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4810_ _7493_/Q _4809_/S _4811_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_2291 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_5790_ _5790_/A1 _5790_/A2 _5791_/A4 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_61_475 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_175_812 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4741_ hold271/Z _4753_/I1 _4741_/S _4741_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XTAP_1590 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_7460_ hold33/Z _7853_/RN _7461_/CLK _7460_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
X_4672_ _7462_/Q _3879_/Z _4672_/B _4673_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_119_238 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_6411_ _6547_/A1 _6417_/A2 _6411_/B _7834_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_174_388 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7391_ _7391_/D _7900_/RN _7767_/CLK _7391_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
X_6342_ hold433/Z _6349_/A2 _6343_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_6273_ _6545_/A1 _6281_/A2 _6273_/B hold105/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_5224_ _5302_/A1 _5195_/B _5224_/A3 _5224_/A4 _5687_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__or4_4
XFILLER_115_499 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_130_469 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_69_542 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5155_ _5774_/A1 _5643_/A2 _5155_/B _5769_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_111_683 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_29_428 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5086_ _5648_/A1 _5087_/B _5682_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_110_193 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_84_534 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4106_ _4106_/A1 _4106_/A2 _4106_/A3 _4106_/A4 _4107_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand4_2
XFILLER_112_25 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_72_729 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4037_ _7551_/Q _4284_/A1 _4038_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_64_280 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_169_105 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_80_740 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_106 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
X_5988_ _5988_/A1 hold5/Z _6004_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_4
XPHY_139 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_128 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_24_166 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_117 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
X_4939_ _4900_/Z _4915_/Z _5199_/B _4973_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi21_4
X_7727_ _7727_/D _7877_/RN _7747_/CLK hold69/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
X_7658_ _7658_/D _7938_/RN _7738_/CLK _7658_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
X_6609_ _6953_/A1 _6609_/A2 _6611_/A2 _6908_/A1 _7914_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai22_1
XFILLER_119_783 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7589_ _7589_/D _7900_/RN _7592_/CLK _7999_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_134_742 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_21_77 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_137_77 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_97_37 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_121_425 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xoutput180 _3694_/ZN mgmt_gpio_oeb[18] VDD VSS gf180mcu_fd_sc_mcu7t5v0__buf_4
Xoutput191 _3684_/ZN mgmt_gpio_oeb[28] VDD VSS gf180mcu_fd_sc_mcu7t5v0__buf_4
XFILLER_75_501 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xclkbuf_leaf_91_csclk _7407_/CLK _7410_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_153_87 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_75_523 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_75_567 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_16_601 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_15_144 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XPHY_8 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_70_261 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_70_250 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_156_344 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_117_709 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_171_303 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_144_517 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_7_354 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xclkbuf_leaf_44_csclk clkbuf_3_7__f_csclk/Z _7601_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_7_398 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_152_550 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_125_764 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_125_753 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_112_403 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_604 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_615 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
Xclkbuf_leaf_59_csclk clkbuf_3_6__f_csclk/Z _7720_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_87_70 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_626 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_637 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_648 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_659 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_140_789 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_87_92 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_66_534 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_66_523 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_38_247 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6960_ _7692_/Q _7194_/A2 _7188_/A2 _7375_/Q _7782_/Q _7202_/B1 _6967_/A1 VDD VSS
+ gf180mcu_fd_sc_mcu7t5v0__aoi222_1
X_5911_ hold64/Z _5919_/A2 hold93/Z hold94/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_6891_ _7408_/Q _6891_/A2 _6891_/B1 _7508_/Q _6891_/C1 _7394_/Q _6895_/A1 VDD VSS
+ gf180mcu_fd_sc_mcu7t5v0__aoi222_1
XFILLER_179_436 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_179_425 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5842_ hold823/Z _5845_/A2 _5843_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_5773_ _5658_/B _5606_/B _5773_/B _5773_/C _5775_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XFILLER_21_136 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_7512_ _7512_/D _7959_/RN _7959_/CLK _7517_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_166_108 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_148_812 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4724_ hold415/Z _4731_/A2 hold416/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_7443_ _7443_/D _7853_/RN _7603_/CLK _7443_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
X_4655_ _3879_/Z hold47/Z _4656_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_107_219 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_162_325 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xinput60 mgmt_gpio_in[31] input60/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XFILLER_128_591 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
Xinput71 mgmt_gpio_in[8] input71/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyb_1
Xinput82 spi_sdoenb _3663_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyb_1
Xhold811 hold811/I _7522_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
Xhold800 _7530_/Q hold800/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
X_7374_ _7374_/D _7875_/RN _7874_/CLK _7374_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
X_4586_ _6539_/A1 _4588_/A2 _4586_/B _7397_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
Xhold844 _7660_/Q hold844/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
X_6325_ hold611/Z _6332_/A2 _6326_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
Xhold822 _7471_/Q hold822/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
Xinput93 trap input93/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
Xhold833 _7402_/Q hold833/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
Xhold855 _7398_/Q hold855/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
XFILLER_131_712 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_130_211 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_103_425 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xhold877 _7775_/Q hold877/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
Xhold888 hold888/I _7524_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
Xhold866 _7406_/Q hold866/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
X_6256_ _6545_/A1 _6264_/A2 _6256_/B hold175/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_107_69 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
Xhold899 hold899/I _4492_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
X_6187_ _4476_/I _6191_/A2 _6187_/B hold228/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_5207_ _5203_/I _5207_/A2 _5392_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_5138_ _4365_/Z _5138_/A2 _5209_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_111_491 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_123_68 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_57_567 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5069_ _4906_/Z _5069_/A2 _5210_/B _5069_/A4 _5458_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand4_4
XFILLER_72_515 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_38_792 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_72_548 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_25_486 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_52_250 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_139_812 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_9_619 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_40_478 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_166_653 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_148_32 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_32_32 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_165_141 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_148_65 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_126_506 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_113_2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_107_775 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_122_734 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_121_277 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_76_810 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_67_309 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_48_534 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_180_41 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_36_707 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_57_73 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_90_389 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_73_83 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_71_570 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_31_412 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_31_434 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_43_283 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_148_108 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_8_663 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_144_336 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4440_ _7901_/RN _4334_/Z _4440_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__and2_1
Xhold107 _5853_/Z _7573_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
XFILLER_171_144 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_144_347 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
Xhold118 hold118/I _7671_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
Xhold129 hold129/I _6200_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
X_4371_ _4922_/A3 _4922_/A4 _4924_/A1 _4924_/A2 _4374_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor4_1
XFILLER_113_712 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6110_ hold922/Z _6123_/A2 hold923/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_112_211 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7090_ _7851_/Q _7193_/A2 _7193_/B1 _7633_/Q _7193_/C1 _7729_/Q _7097_/A1 VDD VSS
+ gf180mcu_fd_sc_mcu7t5v0__aoi222_1
XTAP_423 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_401 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_412 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_6041_ _6539_/A1 _6055_/A2 _6041_/B _7660_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_85_106 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_456 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_467 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_445 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_434 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_489 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_478 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_27_707 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_39_567 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7992_ _7992_/I _7992_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_94_673 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_66_386 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_54_515 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6943_ _7194_/A2 _7189_/B1 _7201_/B1 _7190_/C1 _6946_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor4_1
XFILLER_34_250 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6874_ _7184_/A1 _6767_/C _7433_/Q _6875_/B2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_5825_ _6545_/A1 _5827_/A2 _5825_/B _7561_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_179_288 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_167_428 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_5756_ _5756_/A1 _5756_/A2 _5756_/A3 _7543_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__or3_1
XFILLER_163_612 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_148_664 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_147_141 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4707_ hold506/Z _4718_/A1 hold507/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_5687_ _5689_/A1 _5689_/A2 _5687_/B _5687_/C _5688_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi211_1
X_7426_ _7426_/D _7923_/RN _7599_/CLK _7983_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
X_4638_ _3830_/Z hold16/Z _4639_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_1
Xhold630 _7718_/Q hold630/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
Xhold663 hold663/I _7714_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
Xhold652 _7670_/Q hold652/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
XFILLER_89_423 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
Xhold641 _7702_/Q hold641/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
XFILLER_78_17 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
Xmax_cap360 input75/Z _7875_/RN VDD VSS gf180mcu_fd_sc_mcu7t5v0__buf_20
X_7357_ _7357_/D _7961_/RN _7570_/CLK _7357_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffsnq_1
X_4569_ _4569_/A1 _6537_/A2 _4573_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
Xhold696 _7872_/Q hold696/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
XFILLER_104_734 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_103_233 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_89_445 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xhold685 _7784_/Q hold685/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
X_6308_ hold423/Z _6315_/A2 _6309_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_7288_ hold803/Z _7289_/A2 _7289_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
Xhold674 hold674/I _7732_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
X_6239_ _7754_/Q hold6/Z _6240_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_134_34 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_131_553 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_103_288 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_990 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_45_526 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_72_356 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_17_239 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_72_389 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_150_99 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_13_434 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_25_283 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_41_721 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_53_570 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_159_53 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_41_798 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_138_141 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_138_174 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_153_144 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_5_633 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_4_176 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_122_531 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_49_810 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_110_737 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_76_673 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_75_150 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_90_120 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3940_ _3940_/A1 _3940_/A2 _3940_/A3 _3940_/A4 _3954_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand4_2
XFILLER_16_250 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_17_773 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_149_428 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3871_ _4212_/A2 hold54/Z _6316_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_4
XFILLER_31_220 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_32_754 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_176_247 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5610_ _5602_/Z _5610_/A2 _5610_/A3 _5609_/Z _5610_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__and4_1
XFILLER_31_286 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6590_ _6590_/A1 _6665_/A2 _6879_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_2
X_5541_ _5369_/B _5024_/Z _5543_/B _5541_/A4 _5550_/C VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor4_2
XFILLER_129_141 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_76_2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_145_623 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_129_174 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5472_ _5668_/A2 _5462_/Z _5472_/B _5472_/C _5474_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi211_1
X_7211_ _7433_/Q _7939_/Q _7211_/B _7213_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_4423_ input85/Z input58/Z _7980_/Q _4423_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_7142_ _7789_/Q _7202_/B1 _7205_/A2 _7739_/Q _7144_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_4354_ _6908_/A1 _7913_/Q _6953_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_4
X_7073_ _7736_/Q _7205_/A2 _7205_/B1 _7744_/Q _7075_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_4285_ _7344_/Q _3734_/Z _4288_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_113_586 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6024_ hold47/Z _6038_/A2 _6024_/B _7652_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_101_759 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_100_247 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_39_353 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_104_37 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_7975_ _7975_/D _7328_/Z _4415_/A2 _7975_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XTAP_2109 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1419 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1408 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_82_676 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6926_ _6937_/A1 _6951_/A2 _7203_/B1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_4
XFILLER_35_570 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_54_389 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6857_ _7527_/Q _6885_/B1 _6890_/A2 _7474_/Q _6859_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_167_247 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6788_ _7803_/Q _6883_/A2 _6883_/B1 _7787_/Q _6791_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_5808_ hold749/Z _5811_/A2 _5809_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_5739_ _5739_/A1 _5739_/A2 _5739_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_13_34 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_10_459 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_129_34 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_108_325 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_13_89 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_135_144 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_150_103 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7409_ _7409_/D _7875_/RN _7410_/CLK _7409_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_150_147 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_145_33 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
Xhold460 hold460/I _7873_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
XFILLER_104_531 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xhold471 hold471/I _4502_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
XFILLER_145_55 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
Xhold493 hold493/I _7598_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
Xhold482 _7585_/Q hold482/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
XFILLER_104_564 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_104_553 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_89_286 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_180_2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_92_418 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_57_161 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_45_367 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_45_378 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1942 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1931 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1920 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_159_737 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1986 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1975 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1964 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1953 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_13_231 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_158_247 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1997 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_146_409 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_13_286 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_139_494 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_127_623 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
Xclkbuf_2_2__f_mgmt_gpio_in[4] clkbuf_0_mgmt_gpio_in[4]/Z _4415_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_181_283 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_126_188 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_5_496 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_79_82 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_79_93 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_150_670 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_110_534 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_96_724 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_95_201 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_4070_ _4284_/A1 _7224_/I0 _4073_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_64_676 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_36_356 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4972_ _5006_/C _5608_/A1 _5714_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_2
X_7760_ _7760_/D _7901_/RN _7858_/CLK _7760_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffsnq_1
XFILLER_17_570 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_36_389 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7691_ _7691_/D _7923_/RN _7698_/CLK _7691_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
X_6711_ _7686_/Q _6884_/B1 _6716_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_3923_ _7828_/Q _6384_/A1 _6418_/A1 _7844_/Q _3943_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_3854_ hold76/I hold54/I _6226_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_4
X_6642_ _6878_/A2 _7909_/Q _7908_/Q _6663_/A4 _6882_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor4_4
XFILLER_177_567 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_177_556 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_165_718 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_149_247 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_158_770 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3785_ hold87/Z _7337_/Q _7414_/Q hold88/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_6573_ _7434_/Q _6633_/A2 _6574_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_5524_ _5524_/I _5558_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_117_144 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_172_250 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_132_103 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5455_ _5648_/A2 _4996_/Z _5643_/A2 _5705_/A2 _5657_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_132_125 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4406_ _7963_/Q _4334_/Z _4407_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_5386_ _5669_/B _5669_/A1 _5292_/B _5621_/B _5716_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_7125_ _7780_/Q _7200_/A2 _7201_/B1 _7674_/Q _7200_/B1 _7868_/Q _7128_/A2 VDD VSS
+ gf180mcu_fd_sc_mcu7t5v0__aoi222_1
X_4337_ _5903_/A2 _4338_/A2 _4438_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_115_36 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_99_595 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_59_415 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_101_567 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_87_779 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_86_245 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7056_ _7001_/C _7933_/Q _7058_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_4268_ _7692_/Q _6107_/A1 _4769_/A1 _7472_/Q _4271_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_6007_ hold47/Z _6021_/A2 _6007_/B _7644_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_27_323 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4199_ _7887_/Q _6520_/A1 _5988_/A1 _7637_/Q _5841_/A1 _7570_/Q _4201_/A1 VDD VSS
+ gf180mcu_fd_sc_mcu7t5v0__aoi222_1
XFILLER_55_643 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_131_46 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1205 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_7958_ _7958_/D _7959_/RN _7959_/CLK _7958_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_131_68 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_82_495 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_82_484 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_82_473 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1238 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1227 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1216 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_152_6 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7889_ _7889_/D _7900_/RN _7897_/CLK _7889_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffsnq_1
XTAP_1249 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_6909_ _6953_/A2 _6941_/A2 _6908_/Z _7194_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor3_4
XFILLER_24_11 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_168_534 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_7_706 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_50_392 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_40_32 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_163_283 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_156_76 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_6_2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_77_212 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xhold290 hold290/I _7828_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
XFILLER_65_73 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_45_153 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_46_676 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_18_389 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1761 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1750 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_60_134 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_60_123 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_45_197 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_1783 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1794 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1772 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_174_504 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_139_291 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_127_420 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_154_250 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_170_743 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_142_412 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_114_125 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5240_ _5385_/B2 _5687_/B _5690_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_2
X_5171_ _5171_/A1 _5171_/A2 _5171_/A3 _5171_/A4 _5191_/B1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand4_1
XFILLER_68_201 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_39_2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_69_779 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4122_ _4141_/A1 _3869_/I _4883_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_4053_ _7761_/Q _6248_/A1 _6384_/A1 _7825_/Q _7841_/Q _6418_/A1 _4057_/A1 VDD VSS
+ gf180mcu_fd_sc_mcu7t5v0__aoi222_1
XFILLER_83_215 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xclkbuf_3_0__f_csclk clkbuf_0_csclk/Z _7407_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
Xinput3 debug_out input3/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XFILLER_49_470 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_64_451 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_36_131 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_52_602 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7812_ _7812_/D _7853_/RN _7812_/CLK _7812_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_64_473 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_52_635 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4955_ _4943_/Z _4955_/A2 _4957_/A4 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_7743_ _7743_/D _7877_/RN _7747_/CLK hold68/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_91_292 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_40_808 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3906_ _3906_/A1 _3906_/A2 _3906_/A3 _3906_/A4 _3917_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand4_1
X_7674_ _7674_/D _7938_/RN _7738_/CLK _7674_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
X_4886_ hold791/Z _4887_/A2 hold792/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_32_392 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_177_386 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3837_ hold38/Z hold89/Z _6022_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_4
X_6625_ _7432_/D _6625_/A2 _6625_/B _7920_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_3768_ hold962/Z _7970_/Q _3772_/S _3768_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_6556_ _7435_/Q _7433_/Q _6556_/B _6557_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_180_529 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_173_570 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5507_ _5648_/A1 _5793_/A2 _5624_/B _5648_/B2 _5649_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_3699_ hold84/I _3699_/ZN VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_105_125 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6487_ hold812/Z _6502_/A2 _6488_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_5438_ _5721_/B _5424_/Z _5438_/A3 _5439_/A4 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor3_1
XFILLER_105_136 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xoutput340 _7503_/Q wb_dat_o[7] VDD VSS gf180mcu_fd_sc_mcu7t5v0__buf_4
X_5369_ _3728_/I _4996_/Z _5369_/B _5370_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_133_489 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_59_212 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_120_139 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_99_392 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7108_ _7433_/Q _7935_/Q _7106_/Z _7108_/B2 _7109_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_7039_ _7035_/Z _7039_/A2 _7039_/A3 _7039_/A4 _7054_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand4_1
XFILLER_142_56 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_142_34 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_19_77 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_19_88 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_83_760 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_83_771 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_28_676 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_43_602 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_82_270 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_35_32 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1002 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1013 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1035 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1046 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_15_337 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_43_668 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1024 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1079 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1068 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1057 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_30_318 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_168_342 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_168_353 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_143_2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_129_707 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_70_498 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_156_526 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_11_565 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_51_86 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_136_250 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_136_283 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_98_808 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_808 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_151_286 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_819 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_105_692 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_76_50 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_38_407 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_65_215 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_46_440 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_46_495 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2270 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_22_808 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2292 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2281 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_4740_ hold865/Z _4740_/I1 _4741_/S _7456_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XTAP_1591 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1580 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_14_381 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_14_392 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4671_ _3879_/Z hold16/Z _4672_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_119_228 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6410_ hold444/Z _6417_/A2 _6411_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_7390_ _7390_/D input75/Z _7410_/CLK _7390_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_162_529 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6341_ _6545_/A1 _6349_/A2 _6341_/B _7801_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_155_570 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_127_283 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_127_294 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6272_ hold104/Z _6281_/A2 _6273_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_5223_ _5302_/A1 _5195_/B _5224_/A3 _5224_/A4 _5433_/C VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor4_4
XFILLER_88_329 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_88_318 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5154_ _5496_/A1 _5543_/B _5153_/C _5552_/A3 _5155_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor4_2
XFILLER_102_128 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_69_554 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4105_ _4105_/A1 _4105_/A2 _4106_/A4 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_5085_ _5496_/A1 _5319_/C _5660_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_110_183 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4036_ _4025_/Z _4036_/A2 _4036_/A3 _4036_/A4 _4036_/ZN VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor4_1
XFILLER_112_37 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_65_771 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_25_657 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_107 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
X_5987_ _6553_/A1 _5987_/A2 _5987_/B _7635_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
XPHY_129 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_12_318 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_40_605 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_118 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
X_4938_ _4941_/C _4941_/B _4942_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_166_802 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7726_ _7726_/D _7853_/RN _7726_/CLK _7726_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffsnq_1
XFILLER_52_498 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_178_673 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_177_161 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7657_ _7657_/D _7923_/RN _7816_/CLK _7657_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
X_4869_ hold398/Z _4872_/A2 hold399/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_6608_ _6586_/B _6608_/A2 _6611_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_118_250 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_7588_ _7588_/D _7900_/RN _7592_/CLK _7998_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_21_34 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6539_ _6539_/A1 _6553_/A2 _6539_/B _7894_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_161_540 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_106_456 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_106_445 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_97_27 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_133_286 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xoutput170 _4433_/Z irq[2] VDD VSS gf180mcu_fd_sc_mcu7t5v0__buf_4
Xoutput181 _3693_/ZN mgmt_gpio_oeb[19] VDD VSS gf180mcu_fd_sc_mcu7t5v0__buf_4
Xoutput192 _3683_/ZN mgmt_gpio_oeb[29] VDD VSS gf180mcu_fd_sc_mcu7t5v0__buf_4
XFILLER_121_448 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_734 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_102_673 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_101_150 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_75_513 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_789 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_47_215 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_63_708 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_62_229 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_43_410 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XPHY_9 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_16_646 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_55_292 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_31_605 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_157_802 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_102_92 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_62_52 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_31_638 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_129_515 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_8_812 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_11_351 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_156_389 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_137_570 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_109_283 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_98_605 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_605 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_616 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_627 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_638 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_649 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_66_546 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_38_237 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_93_354 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5910_ hold92/Z _5919_/A2 hold93/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_34_410 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_53_207 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6890_ _7475_/Q _6890_/A2 _6890_/B1 _7396_/Q _6896_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_46_270 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5841_ _5841_/A1 _6537_/A2 _5845_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_22_605 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5772_ _5772_/A1 _5173_/B _5772_/A3 _5773_/C VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_34_498 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7511_ _7511_/D _7959_/RN _7959_/CLK _7511_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffsnq_1
X_4723_ _4454_/Z _4731_/A2 _4723_/B _7445_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_7442_ _7442_/D _7853_/RN _7603_/CLK _7442_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_30_682 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4654_ hold514/Z _4685_/A1 hold515/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_175_698 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
Xinput61 mgmt_gpio_in[32] input61/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyb_1
Xinput50 mgmt_gpio_in[22] input50/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyb_1
Xinput72 mgmt_gpio_in[9] input72/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyc_1
Xhold812 _7870_/Q hold812/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
Xhold801 hold801/I _4877_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
X_7373_ _7373_/D _7875_/RN _7822_/CLK _7373_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
X_4585_ hold769/Z _4588_/A2 _4586_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_143_540 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6324_ _6545_/A1 _6332_/A2 _6324_/B hold166/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
Xinput83 spimemio_flash_clk input83/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyb_1
Xhold823 _7569_/Q hold823/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
Xinput94 uart_enabled _4400_/S VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyb_1
Xhold834 _7477_/Q hold834/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
Xhold845 _7766_/Q hold845/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
X_6255_ hold173/Z _6264_/A2 hold174/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_107_37 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_89_638 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xhold856 _7372_/Q hold856/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
Xhold889 _7469_/Q hold889/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
Xhold867 _7547_/Q hold867/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
Xhold878 _7759_/Q hold878/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
XFILLER_170_392 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5206_ _5369_/B _5206_/A2 _5205_/Z _5207_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor3_1
XFILLER_115_286 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_67_19 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6186_ hold227/Z _6191_/A2 _6187_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_131_779 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5137_ _5309_/A1 _3723_/I _5344_/A1 _5498_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand3_4
XFILLER_84_321 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_29_215 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_57_524 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5068_ _5302_/A1 _5211_/A3 _4920_/Z _5069_/A4 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_123_47 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_57_579 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_84_398 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4019_ _7656_/Q _6022_/A1 _5971_/A1 _7632_/Q _4020_/A4 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_16_34 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_25_410 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_25_476 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_40_402 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_52_262 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_40_424 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7709_ _7709_/D _7877_/RN _7722_/CLK _7709_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffsnq_1
XFILLER_8_108 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_21_682 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_166_676 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_154_805 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_180_112 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_138_389 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_119_570 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_106_2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_107_798 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_164_54 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_121_212 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_79_148 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_76_800 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_87_170 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_597 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_75_354 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_75_332 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_90_302 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_63_538 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_35_229 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_113_80 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_73_73 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_16_454 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_129_312 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_172_602 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_156_142 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_7_141 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xhold108 _7667_/Q hold108/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
X_4370_ _4924_/A3 _4924_/A4 _4370_/A3 _4370_/A4 _4372_/A4 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor4_1
XFILLER_125_540 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
Xhold119 _7651_/Q hold119/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
XFILLER_152_392 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_152_381 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_98_424 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_424 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_402 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_413 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_6040_ hold844/Z _6055_/A2 _6041_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_79_660 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_67_811 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_457 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_446 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_435 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_94_630 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_66_321 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_479 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_468 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_21_2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7991_ _7991_/I _7991_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_6942_ _7189_/A2 _7191_/A2 _7197_/A2 _7193_/B1 _6946_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor4_1
XFILLER_19_281 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_179_212 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_81_357 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6873_ _6873_/A1 _6867_/Z _6873_/A3 _6875_/B1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_50_700 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5824_ hold157/Z _5827_/A2 _5825_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_22_402 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_50_744 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_139_109 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5755_ _5755_/A1 _5755_/A2 _5777_/B _5756_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi21_1
Xclkbuf_leaf_90_csclk _7407_/CLK _7570_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_148_676 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4706_ _4718_/A1 _4706_/A2 _4706_/B hold322/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_5686_ _5363_/B _5686_/A2 _5627_/Z _5686_/A4 _5686_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__and4_1
XFILLER_147_164 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4637_ hold483/Z _4652_/A1 hold484/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_7425_ _7425_/D _7853_/RN _7818_/CLK _7425_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_163_668 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_162_123 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_151_808 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xhold620 _7684_/Q hold620/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
XFILLER_150_318 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_104_724 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
Xhold653 _7654_/Q hold653/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
Xhold642 hold642/I _6130_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
X_7356_ _7356_/D input75/Z _7570_/CLK _7356_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffsnq_1
Xhold631 _7365_/Q hold631/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
X_4568_ _4454_/Z _4568_/A2 _4568_/B _7390_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_103_223 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_103_212 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xhold675 _7768_/Q hold675/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
Xhold686 _7824_/Q hold686/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
X_6307_ _6545_/A1 _6315_/A2 _6307_/B hold103/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
Xhold697 _8003_/I hold697/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
Xhold664 _7876_/Q hold664/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
X_7287_ hold47/Z _7289_/A2 _7287_/B _7960_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_4499_ hold745/Z _4504_/A2 hold746/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_6238_ _4476_/I hold6/Z _6238_/B hold218/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_77_608 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6169_ hold348/Z _6174_/A2 _6170_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_980 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_85_641 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_991 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_57_354 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_84_173 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_72_313 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_57_376 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_150_34 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xclkbuf_leaf_43_csclk clkbuf_3_7__f_csclk/Z _7821_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_60_508 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_40_210 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_13_457 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_13_446 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
Xclkbuf_leaf_58_csclk clkbuf_3_6__f_csclk/Z _7816_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_9_428 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_40_254 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_154_602 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_138_120 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_166_473 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_153_101 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_181_454 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_181_432 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_142_808 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_141_307 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_134_392 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_4_37 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_68_62 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_110_727 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_48_310 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_383 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_48_321 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_48_387 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_36_538 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_84_94 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_63_357 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_90_176 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3870_ _4075_/B _3869_/I _4505_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_4
XFILLER_32_744 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_290 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
X_5540_ _5735_/A2 _5179_/B _5540_/B1 _5540_/B2 _5540_/C _5642_/A4 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi221_2
X_5471_ _5674_/A1 _5471_/A2 _5749_/A3 _5471_/A4 _5472_/C VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand4_1
XFILLER_69_2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4422_ _4422_/I _4422_/ZN VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_7210_ _7210_/A1 _7210_/A2 _7210_/B _7433_/Q _7211_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XFILLER_160_605 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_132_318 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7141_ _7877_/Q _7195_/C1 _7193_/C1 _7731_/Q _7667_/Q _7194_/B1 _7144_/A2 VDD VSS
+ gf180mcu_fd_sc_mcu7t5v0__aoi222_1
X_4353_ _6905_/A1 _7916_/Q _6937_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_4
X_7072_ _7826_/Q _7202_/A2 _7204_/B1 _7770_/Q _7077_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_4284_ _4284_/A1 _4427_/B _7219_/A1 _4284_/B _7548_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai31_1
X_6023_ hold691/Z _6038_/A2 _6024_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_100_259 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_67_641 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_94_460 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7974_ _7974_/D _7327_/Z _4415_/A2 _7974_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XTAP_1409 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_81_154 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6925_ _7912_/Q _7911_/Q _6936_/A2 _6951_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand3_4
XFILLER_120_37 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_35_560 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_80_19 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6856_ _7529_/Q _6881_/A2 _6881_/B1 _7523_/Q _6859_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_167_226 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_167_215 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6787_ _6787_/A1 _6787_/A2 _6787_/A3 _6792_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand3_1
X_3999_ _3999_/A1 _3999_/A2 _3999_/A3 _3998_/Z _7227_/I0 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand4_4
X_5807_ _5807_/A1 _6537_/A2 _5811_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_148_451 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5738_ _5698_/B _5738_/A2 _5738_/B _5738_/C _5756_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_136_646 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5669_ _5669_/A1 _5179_/B _5669_/B _5799_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_7408_ _7408_/D input75/Z _7637_/CLK _7408_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
X_7339_ _7339_/D _7294_/Z _7972_/CLK _7339_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_151_638 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_150_115 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
Xhold461 _7825_/Q hold461/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
XFILLER_116_392 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_89_221 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xhold450 hold450/I _6394_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
Xhold472 hold472/I _7361_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
Xhold494 _7708_/Q hold494/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
Xhold483 _7994_/I hold483/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
XFILLER_161_55 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_173_2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_72_110 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_18_549 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_1910 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_45_357 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1943 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1932 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1921 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_72_187 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_72_176 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1976 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1965 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1954 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_14_744 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1998 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1987 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_14_788 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_41_574 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_110_81 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_70_52 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_126_101 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_70_63 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_154_421 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_142_605 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_107_392 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_96_747 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_95_224 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_68_427 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_49_641 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_95_268 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_76_471 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_76_460 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_48_162 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_64_622 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_64_666 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4971_ _5006_/B _5254_/A2 _5206_/A2 _5104_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor3_4
XFILLER_91_496 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6710_ _7133_/S _6710_/A2 _6710_/B _7922_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_7690_ _7690_/D _7923_/RN _7815_/CLK _7690_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_32_530 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3922_ _4402_/A1 _4427_/B _3922_/B hold945/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_149_226 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_149_237 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_149_215 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3853_ _4212_/A2 hold82/Z _6452_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_4
X_6641_ _7910_/Q _6663_/A4 _6658_/A3 _6885_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor3_4
XFILLER_20_747 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3784_ _3810_/S _3781_/Z hold25/Z hold26/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi21_4
XFILLER_118_602 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6572_ _6572_/A1 _4352_/B _6618_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_2
X_5523_ _5519_/B _5559_/A1 _5523_/A3 _5524_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__or3_1
X_5454_ _5783_/A2 _5668_/A2 _5454_/B _5460_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_133_627 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_132_137 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5385_ _5603_/A1 _4993_/B _4993_/C _5409_/B2 _5385_/B2 _5583_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai32_1
X_4405_ _7424_/Q input3/Z input1/Z _4405_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_4336_ _7978_/Q hold21/I _4338_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_87_703 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_7124_ _7884_/Q _7203_/B1 _7204_/A2 _7844_/Q _7129_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_141_682 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_59_405 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_7055_ _7607_/Q _7210_/A2 _7055_/B _7433_/Q _7058_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi211_1
X_4267_ _4267_/A1 _4267_/A2 _4267_/A3 _4267_/A4 _4281_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand4_1
X_6006_ hold584/Z _6021_/A2 _6007_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_4198_ _4198_/A1 _4198_/A2 _4198_/A3 _4198_/A4 _4202_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand4_1
XFILLER_55_600 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_67_482 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_67_493 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_39_195 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_82_463 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_27_357 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7957_ _7957_/D _7959_/RN _7959_/CLK _7957_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XTAP_1239 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1228 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1217 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1206 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_70_636 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_54_176 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7888_ _7888_/D _7900_/RN _7896_/CLK _7888_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
X_6908_ _6908_/A1 _7913_/Q _6908_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__or2_4
XFILLER_168_513 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_168_524 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6839_ _6839_/A1 _6839_/A2 _6839_/A3 _6848_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_176_590 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_156_33 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_136_465 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_124_605 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_108_156 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_156_88 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_108_189 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_2_412 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_156_99 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xhold280 _7884_/Q hold280/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
Xhold291 _7772_/Q hold291/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
XFILLER_78_747 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_77_235 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_65_419 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_58_460 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_105_70 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_18_346 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_73_496 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_33_327 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1751 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1740 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_61_658 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_14_530 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1784 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1773 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1762 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_60_179 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1795 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_81_73 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_81_84 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_41_371 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_154_273 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_115_649 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_115_638 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_114_104 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_69_703 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_5_283 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_170_788 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_5170_ _5666_/A1 _5658_/B _5179_/B _5672_/A2 _5171_/A4 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_69_714 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_122_192 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_110_321 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_96_555 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_96_544 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4121_ hold82/Z _3959_/Z _4589_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_4052_ _4052_/A1 _4052_/A2 _4052_/A3 _4058_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_84_717 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_77_780 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xinput4 mask_rev_in[0] input4/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XFILLER_49_482 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_7811_ _7811_/D _7853_/RN _7811_/CLK _7811_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_64_463 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_36_176 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_51_102 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4954_ _5069_/A2 _4930_/Z _4953_/Z _5661_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand3_4
X_7742_ _7742_/D _7877_/RN _7872_/CLK _7742_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffsnq_1
X_3905_ input60/Z _5886_/A1 _6537_/A1 _7901_/Q _3906_/A4 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_177_354 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7673_ _7673_/D _7923_/RN _7698_/CLK _7673_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
X_4885_ hold47/Z _4887_/A2 _4885_/B hold407/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_20_522 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_32_382 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6624_ _7920_/Q _6625_/A2 _6625_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_3836_ hold38/Z hold42/Z _5937_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_4
X_3767_ _7970_/Q hold960/Z _3772_/S _3767_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_20_588 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6555_ _7435_/Q _7433_/Q _6562_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_5506_ _5735_/A2 _5179_/B _5540_/C _5506_/C _5508_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XFILLER_106_605 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_160_210 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_145_262 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3698_ _7719_/Q _3698_/ZN VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_6486_ _6486_/A1 _6537_/A2 _6502_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_4
X_5437_ _5714_/B1 _5722_/A1 _5437_/B _5438_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
Xoutput330 _7945_/Q wb_dat_o[27] VDD VSS gf180mcu_fd_sc_mcu7t5v0__buf_4
Xoutput341 _7486_/Q wb_dat_o[8] VDD VSS gf180mcu_fd_sc_mcu7t5v0__buf_4
X_5368_ _5689_/A1 _5618_/B1 _5565_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_4319_ _4309_/S _4319_/A2 _4319_/B _7338_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_5299_ _5173_/C _5299_/A2 _5299_/A3 _5299_/A4 _5300_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand4_1
XFILLER_113_170 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7107_ _7107_/A1 _7210_/A2 _7433_/Q _7108_/B2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_7038_ _7817_/Q _7207_/A2 _7205_/B1 hold68/I _7039_/A4 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_101_354 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_74_205 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_75_739 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_142_79 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_67_290 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_28_666 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_83_783 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_27_176 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1003 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_169_800 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_1036 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1047 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1014 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1025 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_168_321 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1069 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1058 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_35_99 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_42_179 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_136_2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_164_560 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_137_774 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_51_98 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_136_262 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_152_744 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_124_457 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_809 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_111_129 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_104_181 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_78_544 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_120_663 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_76_62 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_59_780 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_81_709 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_74_761 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_61_400 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_18_176 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_46_463 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2271 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2260 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_18_198 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_2293 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2282 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_92_94 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_159_354 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1592 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1581 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1570 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_61_499 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_147_516 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4670_ hold381/Z _4685_/A1 hold382/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_128_763 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6340_ hold169/Z _6349_/A2 _6341_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_51_2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_143_766 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_6271_ _4460_/Z _6281_/A2 _6271_/B _7768_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_6_592 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5222_ _5376_/B _5392_/B2 _5294_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_115_479 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_102_118 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_69_511 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5153_ _5552_/A3 _5539_/A3 _5543_/B _5153_/C _5180_/C1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XFILLER_123_490 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_111_641 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4104_ _4104_/A1 _4104_/A2 _4104_/A3 _4104_/A4 _4105_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand4_1
XFILLER_69_566 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5084_ _5643_/A2 _5087_/B _5600_/B2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_110_195 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4035_ _4035_/A1 _4035_/A2 _4035_/A3 _4035_/A4 _4036_/A4 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand4_1
XFILLER_65_783 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_64_260 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_80_731 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_25_647 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_37_496 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5986_ hold312/Z _5987_/A2 _5987_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XPHY_119 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_108 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
X_4937_ _5200_/B _3727_/I _4946_/A1 _5230_/A1 _4941_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor4_4
X_7725_ _7725_/D _7877_/RN _7747_/CLK _7725_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffsnq_1
XFILLER_24_179 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_177_140 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7656_ _7656_/D _7923_/RN _7736_/CLK _7656_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_20_341 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4868_ _4868_/A1 _7285_/A2 _4872_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_3819_ hold609/Z hold27/Z _3819_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__or2_4
X_6607_ _7434_/Q _6610_/A3 _6608_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_165_357 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7587_ _7587_/D _7875_/RN _7874_/CLK _7587_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
X_4799_ _7486_/Q _4809_/S _4800_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_21_79 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6538_ hold788/Z _6553_/A2 _6539_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_137_68 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_134_744 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6469_ _6469_/A1 hold5/Z _6485_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_4
XFILLER_97_17 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_702 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xoutput171 _4409_/ZN mgmt_gpio_oeb[0] VDD VSS gf180mcu_fd_sc_mcu7t5v0__buf_4
Xoutput182 _4407_/ZN mgmt_gpio_oeb[1] VDD VSS gf180mcu_fd_sc_mcu7t5v0__buf_4
Xoutput193 _3710_/ZN mgmt_gpio_oeb[2] VDD VSS gf180mcu_fd_sc_mcu7t5v0__buf_4
XFILLER_87_352 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_768 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_28_463 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_16_658 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_15_168 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_169_641 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_62_64 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_30_105 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_43_499 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_168_140 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_7_312 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_171_316 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_124_276 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_606 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_140_747 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_87_50 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_617 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_628 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_639 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_120_460 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_47_783 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_19_496 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_34_422 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_61_230 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5840_ _6549_/A1 _5840_/A2 _5840_/B _7568_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
XTAP_2090 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_5771_ _5771_/A1 _5805_/A1 _5805_/B _5787_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_99_2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_175_611 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4722_ hold846/Z _4731_/A2 _4723_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_7510_ _7510_/D _7938_/RN _7532_/CLK _7510_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_175_633 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_175_622 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7441_ _7441_/D _7853_/RN _7600_/CLK _7441_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_30_672 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_163_806 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_147_357 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4653_ _4653_/A1 _5903_/A2 _4686_/B1 _3879_/Z hold22/Z _4685_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi221_4
Xinput40 mgmt_gpio_in[13] input40/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XFILLER_174_176 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xinput62 mgmt_gpio_in[33] input62/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XFILLER_128_582 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_116_722 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
Xinput51 mgmt_gpio_in[23] input51/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyb_1
Xinput73 pad_flash_io0_di input73/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyb_1
Xhold802 hold802/I _7530_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
X_7372_ _7372_/D _7875_/RN _7410_/CLK _7372_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
X_4584_ _4584_/A1 _6537_/A2 _4588_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
Xinput95 wb_adr_i[0] _3723_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__buf_16
X_6323_ hold164/Z _6332_/A2 hold165/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
Xinput84 spimemio_flash_csb input84/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyb_1
Xhold813 _7495_/Q hold813/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
Xhold846 _7445_/Q hold846/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
Xhold824 _7508_/Q hold824/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
Xhold835 _7887_/Q hold835/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
XFILLER_143_552 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_107_27 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_88_105 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6254_ _4460_/Z _6264_/A2 _6254_/B _7760_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
Xhold879 _7855_/Q hold879/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
Xhold857 _7390_/Q hold857/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
Xhold868 _7475_/Q hold868/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
X_5205_ _5338_/A1 _4996_/Z _5205_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_103_449 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_103_438 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6185_ hold16/Z _6191_/A2 _6185_/B hold29/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_5136_ _5136_/A1 _5344_/A2 _5680_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_2
XFILLER_97_683 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5067_ _3722_/I _5087_/C _5344_/A1 _5527_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand3_4
XFILLER_45_709 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4018_ input24/Z _4239_/A2 _6282_/A1 _7778_/Q _4020_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_72_528 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_44_208 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_53_731 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_80_583 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_12_105 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5969_ hold139/Z _5970_/A2 _5970_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_25_499 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7708_ _7708_/D _7853_/RN _7722_/CLK _7708_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffsnq_1
XFILLER_32_34 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_148_34 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7639_ _7639_/D _7961_/RN _7639_/CLK _7639_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_165_176 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_148_78 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_181_658 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_107_733 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_180_179 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_164_33 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_122_747 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_94_108 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_102_460 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_76_812 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_57_75 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_90_314 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_29_783 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_35_219 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_43_241 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_31_425 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_31_469 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_169_493 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_145_806 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_129_357 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_172_614 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_156_176 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_8_676 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_7_153 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_172_658 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_171_146 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_144_338 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xhold109 hold109/I _7667_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
XFILLER_113_703 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_403 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_414 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_458 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_447 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_436 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_425 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_121_780 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_469 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_14_2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_27_709 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_39_558 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7990_ _7990_/I _7990_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_93_141 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6941_ _6941_/A1 _6941_/A2 _7196_/B1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_4
XFILLER_62_550 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6872_ _7525_/Q _6889_/A2 _6853_/Z _6830_/B _6872_/C _6873_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi221_1
X_5823_ _4460_/Z _5827_/A2 _5823_/B _7560_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_179_268 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_22_458 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5754_ _5754_/A1 _5754_/A2 _5754_/A3 _5800_/A1 _5755_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor4_1
X_4705_ hold18/Z _3819_/Z _4705_/B _4706_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_5685_ _5759_/A1 _5724_/A2 _5685_/B _5686_/A4 VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_175_496 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4636_ _4652_/A1 hold468/Z _4636_/B hold469/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_7424_ _7424_/D _7853_/RN _7601_/CLK _7424_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_147_176 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_118_37 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
Xhold621 hold621/I _6092_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
X_7355_ _7355_/D input75/Z _7570_/CLK _7355_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffsnq_1
Xhold610 _7606_/Q hold610/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
XFILLER_162_179 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
Xmax_cap351 hold5/Z _7285_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__buf_20
Xhold643 hold643/I _7702_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
XFILLER_89_403 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
Xhold654 _7686_/Q hold654/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
X_6306_ hold102/Z _6315_/A2 _6307_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
Xhold632 hold632/I _4511_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
X_4567_ hold857/Z _4568_/A2 _4568_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
Xhold687 _7630_/Q hold687/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
XFILLER_131_511 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_104_747 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_89_425 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7286_ hold391/Z _7289_/A2 _7287_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_4498_ _6547_/A1 _4504_/A2 _4498_/B hold519/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
Xhold676 _7668_/Q hold676/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
Xhold665 _7814_/Q hold665/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
X_6237_ _7753_/Q hold6/Z _6238_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
Xhold698 _7625_/Q hold698/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
XFILLER_134_58 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6168_ _6547_/A1 _6174_/A2 _6168_/B _7720_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_76_108 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_970 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_5119_ _5476_/B _5689_/A2 _7520_/Q _5519_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
XTAP_981 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_992 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_6099_ hold536/Z _6106_/A2 hold537/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_17_208 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_175_6 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_150_46 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_84_185 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_25_241 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_26_742 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_13_425 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_41_712 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_41_723 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_179_780 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_139_611 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_40_299 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_166_463 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_138_176 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_154_658 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_138_198 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_153_179 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_107_574 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_4_134 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_181_499 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_107_596 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_108_81 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_110_717 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_103_780 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_95_428 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_49_812 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_31_200 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_140_90 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_31_211 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_291 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_280 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_144_102 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5470_ _4969_/C _4996_/Z _5471_/A4 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_172_422 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_157_496 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4421_ _4424_/A1 input86/Z _4422_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_144_179 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_99_712 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7140_ _7140_/A1 _7140_/A2 _7140_/A3 _7140_/A4 _7140_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__and4_1
XFILLER_98_200 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4352_ _7001_/C _4361_/A2 _4352_/B _7433_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_7071_ _7762_/Q _7202_/C2 _7202_/B1 _7786_/Q _7077_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_4283_ _4283_/A1 _4283_/A2 _4283_/A3 _4283_/A4 _7219_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor4_4
X_6022_ _6022_/A1 _7285_/A2 _6038_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_4
XFILLER_58_108 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7973_ _7973_/D _7326_/Z _4415_/A2 _7973_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_66_174 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_81_144 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6924_ _7912_/Q _7911_/Q _6955_/A4 _6908_/Z _7190_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor4_4
XFILLER_23_712 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_168_717 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_62_380 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_6855_ _7531_/Q _6892_/B1 _6880_/B1 _7409_/Q _6867_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_50_531 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6786_ _7697_/Q _6881_/B1 _6880_/B1 _7811_/Q _6787_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_5806_ _5806_/A1 _5806_/A2 _5806_/A3 _5806_/A4 _7545_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand4_1
X_3998_ _3998_/A1 _3998_/A2 _3998_/A3 _3998_/A4 _3998_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__and4_1
X_5737_ _5795_/A2 _5737_/A2 _5785_/A1 _5737_/B _5738_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai31_1
XFILLER_163_400 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_148_463 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5668_ _5783_/A2 _5668_/A2 _5668_/B _5668_/C _5776_/A4 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi211_2
X_7407_ _7407_/D input75/Z _7407_/CLK _7407_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
X_5599_ _5599_/A1 _5661_/B _5656_/A2 _5665_/A1 _5599_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__and4_1
XFILLER_135_168 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4619_ _5886_/A1 _5903_/A2 _4686_/B1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_4
XFILLER_2_605 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7338_ _7338_/D _7293_/Z _7972_/CLK hold87/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_163_499 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_163_488 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_150_105 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xhold462 hold462/I _6392_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
Xhold451 hold451/I _7826_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
Xhold440 hold440/I _7890_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
X_7269_ _7519_/Q _7269_/A2 _7271_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_150_149 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xhold495 hold495/I _6143_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
Xhold484 hold484/I _4640_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
Xhold473 _7369_/Q hold473/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
XFILLER_1_148 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_77_428 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_161_12 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_85_461 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_57_152 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_57_141 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_45_325 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_166_2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1900 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_61_807 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1933 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1922 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1911 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_159_728 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1977 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1966 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1955 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1944 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_159_739 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1999 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1988 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_9_215 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_139_430 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_167_783 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_181_230 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_166_282 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_139_496 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_5_421 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_5_410 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_5_465 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_182_797 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_126_179 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_122_330 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_79_73 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_150_683 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_1_682 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_110_569 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_48_174 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_63_144 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_4970_ _5006_/B _5206_/A2 _5608_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_4
X_3921_ _7554_/Q _4284_/A1 _3921_/B _4427_/B _3922_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XFILLER_44_380 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3852_ hold72/I _4075_/B _4239_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_4
X_6640_ _7910_/Q _6658_/A2 _6662_/A3 _6889_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor3_4
XFILLER_165_709 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_81_2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6571_ _6557_/I _6571_/A2 _6570_/Z _6564_/B _6571_/B2 _7905_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai32_1
X_5522_ _5522_/A1 _5520_/C _5522_/B1 _5522_/B2 _7540_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_3783_ hold24/Z hold193/Z _3810_/S _3783_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_4
XFILLER_173_753 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_5453_ _5714_/A1 _5527_/A1 _5668_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_2
XFILLER_106_809 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5384_ _5392_/A1 _5392_/A2 _5376_/B _5405_/B _5392_/B2 _5702_/C VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai32_1
XFILLER_145_499 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xclkbuf_leaf_42_csclk clkbuf_3_7__f_csclk/Z _7722_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_132_105 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4404_ _7979_/Q _4425_/A2 _4404_/B _4404_/ZN VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_99_531 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4335_ _7630_/Q _4335_/A2 _5903_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_4
X_7123_ _7836_/Q _7203_/A2 _7204_/B1 _7772_/Q _7129_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_5_70 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_113_374 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_101_503 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_59_428 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7054_ _7054_/A1 _7054_/A2 _7054_/A3 _7054_/A4 _7055_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__or4_1
XFILLER_87_759 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_86_247 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4266_ _7830_/Q _6401_/A1 _4614_/A1 _7409_/Q _4267_/A4 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_1
Xclkbuf_leaf_57_csclk clkbuf_3_6__f_csclk/Z _7737_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_67_461 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_6005_ _6005_/A1 _7285_/A2 _6021_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_4
XFILLER_39_141 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4197_ _7895_/Q _6537_/A1 _4594_/A1 _7402_/Q _6243_/A1 _7757_/Q _4198_/A4 VDD VSS
+ gf180mcu_fd_sc_mcu7t5v0__aoi222_1
XFILLER_82_442 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7956_ _7956_/D _7959_/RN _7959_/CLK _7956_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_91_19 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_1229 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1218 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1207 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_6907_ _6953_/A1 _6599_/Z _6941_/A2 _7195_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor3_4
X_7887_ _7887_/D _7900_/RN _7887_/CLK _7887_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
X_6838_ _7382_/Q _6882_/A2 _6882_/B1 _7659_/Q _6839_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_50_383 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_149_783 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_6769_ _7680_/Q _6887_/B1 _6891_/B1 _7672_/Q _6771_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_10_247 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_164_742 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_40_34 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_136_455 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_151_436 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_151_425 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_108_179 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xhold270 hold270/I _7901_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
XFILLER_120_812 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xhold292 hold292/I _7772_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
Xhold281 hold281/I _6517_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
XFILLER_93_707 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_86_770 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_1_17 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_18_325 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_45_144 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_73_486 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_65_97 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1752 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1741 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1730 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_121_70 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_60_125 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1785 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1774 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1763 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1796 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_41_361 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_182_594 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_127_499 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_111_812 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_69_726 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_110_311 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_96_534 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_68_247 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4120_ _4141_/A1 _3881_/Z _4863_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_4051_ _7857_/Q _6452_/A1 _6401_/A1 _7833_/Q _7809_/Q _6350_/A1 _4052_/A3 VDD VSS
+ gf180mcu_fd_sc_mcu7t5v0__aoi222_1
XFILLER_83_239 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xinput5 mask_rev_in[10] input5/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XFILLER_49_472 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7810_ _7810_/D _7853_/RN _7812_/CLK _7810_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_92_795 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_24_317 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4953_ _4906_/Z _5138_/A2 _4953_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__and2_4
XFILLER_91_283 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7741_ _7741_/D _7938_/RN _7741_/CLK _7741_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffsnq_1
XFILLER_178_812 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3904_ input51/Z _4275_/A2 _6469_/A1 _7869_/Q _3906_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_7672_ _7672_/D _7923_/RN _7816_/CLK _7672_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
X_4884_ hold405/Z _4887_/A2 hold406/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_6623_ _7432_/Q _7435_/Q _6623_/B _6625_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_177_388 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3835_ _3783_/Z hold41/Z hold75/I hold71/I hold42/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__or4_4
XFILLER_20_534 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3766_ _7971_/Q hold957/Z _3772_/S _3766_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_6554_ _7433_/Q _4331_/Z _6556_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_5505_ _5155_/B _5505_/A2 _5499_/Z _5505_/A4 _5505_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__or4_1
XFILLER_146_764 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_6485_ _6553_/A1 _6485_/A2 _6485_/B hold241/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_161_712 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_160_200 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3697_ hold69/I _3697_/ZN VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_133_425 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5436_ _5731_/B _5287_/B _5439_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_10_37 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_133_469 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_126_37 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_105_127 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xoutput331 _7946_/Q wb_dat_o[28] VDD VSS gf180mcu_fd_sc_mcu7t5v0__buf_4
Xoutput342 _7487_/Q wb_dat_o[9] VDD VSS gf180mcu_fd_sc_mcu7t5v0__buf_4
Xoutput320 _7480_/Q wb_dat_o[18] VDD VSS gf180mcu_fd_sc_mcu7t5v0__buf_4
X_5367_ _5774_/A1 _5669_/A1 _5782_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_126_48 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_120_108 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_114_672 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_102_812 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_86_19 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_59_203 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4318_ _7337_/Q _7414_/Q _4318_/B _4319_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_141_480 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7106_ _7210_/A2 _7106_/A2 _7106_/A3 _7106_/A4 _7106_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__or4_1
X_5298_ _5580_/A1 _5298_/A2 _5298_/A3 _5298_/A4 _5299_/A4 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor4_2
X_7037_ _7679_/Q _7191_/A2 _7194_/B1 hold79/I _7039_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_87_589 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_87_567 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_75_729 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_19_35 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4249_ input4/Z _4249_/A2 _4764_/A1 _7470_/Q _4253_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_19_79 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_27_144 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_28_656 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_82_250 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_82_261 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1004 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1037 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_7939_ _7939_/D _7961_/RN _7940_/CLK _7939_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XTAP_1015 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1026 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_169_812 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_70_456 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1059 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1048 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_35_89 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_143_4 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_129_709 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_11_567 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_51_33 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_129_2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_109_499 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_3_700 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_3_755 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_105_650 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_104_160 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_78_534 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_2_276 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_76_52 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_78_589 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_74_751 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_19_634 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_19_689 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_2261 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2250 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_132_91 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_73_283 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_178_108 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2294 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2283 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2272 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1560 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1593 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1582 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1571 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_128_742 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_143_712 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_142_200 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_115_425 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_170_531 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_142_211 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6270_ hold675/Z _6281_/A2 _6271_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_5221_ _5585_/A1 _5421_/A1 _5203_/I _5392_/B2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand3_2
XFILLER_102_108 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_44_2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5152_ _5528_/A2 _5020_/Z _5122_/Z _5150_/Z _5546_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand4_2
X_4103_ _7872_/Q _6486_/A1 _6299_/A1 _7784_/Q _6265_/A1 _7768_/Q _4104_/A4 VDD VSS
+ gf180mcu_fd_sc_mcu7t5v0__aoi222_1
X_5083_ _5087_/B _5779_/A1 _5692_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_110_185 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4034_ hold59/I _6435_/A1 _5988_/A1 _7640_/Q _5870_/A1 _7575_/Q _4035_/A4 VDD VSS
+ gf180mcu_fd_sc_mcu7t5v0__aoi222_1
XFILLER_64_250 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5985_ _4481_/I _5987_/A2 _5985_/B _7634_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_7724_ _7724_/D _7877_/RN _7729_/CLK _7724_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffsnq_1
XFILLER_52_478 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_52_467 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_109 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
X_4936_ _5199_/B _5201_/B _4915_/Z _5385_/B2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_33_692 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_178_664 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7655_ _7655_/D _7923_/RN _7735_/CLK _7655_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_20_331 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4867_ _4454_/Z _4867_/A2 _4867_/B hold893/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_3818_ hold609/Z hold27/Z _5903_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_4
XFILLER_119_720 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6606_ _6953_/A2 _6950_/A2 _6610_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_7586_ _7586_/D _7875_/RN _7874_/CLK _7586_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
X_4798_ _7513_/Q _7959_/RN _4809_/S VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_4
X_6537_ _6537_/A1 _6537_/A2 _6553_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_4
XFILLER_20_386 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3749_ input58/Z _7976_/Q _3749_/S _7976_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_134_756 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_134_734 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_6468_ _6553_/A1 _6468_/A2 _6468_/B hold244/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_161_564 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_133_244 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6399_ hold260/Z _6400_/A2 hold261/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_5419_ _5087_/B _5292_/B _5419_/B _5419_/C _5727_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi211_2
Xoutput194 _3682_/ZN mgmt_gpio_oeb[30] VDD VSS gf180mcu_fd_sc_mcu7t5v0__buf_4
XFILLER_121_428 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
Xoutput172 _3702_/ZN mgmt_gpio_oeb[10] VDD VSS gf180mcu_fd_sc_mcu7t5v0__buf_4
Xoutput183 _3692_/ZN mgmt_gpio_oeb[20] VDD VSS gf180mcu_fd_sc_mcu7t5v0__buf_4
XFILLER_102_631 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_101_130 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_153_68 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_101_174 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_47_217 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_47_239 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_83_570 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_71_721 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_55_283 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_169_620 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_71_798 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_70_275 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_178_65 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_7_357 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_125_712 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_152_531 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_152_520 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_124_211 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_124_266 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_112_417 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_3_563 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_607 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_97_128 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_618 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_629 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_94_802 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_87_73 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_93_312 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_39_729 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_19_420 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_19_453 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_46_250 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_62_743 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_179_428 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2091 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2080 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_5770_ _5770_/I _5805_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_61_286 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_159_141 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1390 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_4721_ _6539_/A1 _4731_/A2 _4721_/B _7444_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_4652_ _4652_/A1 _4652_/A2 _4652_/B hold325/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_7440_ _7440_/D _7923_/RN _7599_/CLK _7989_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
Xinput30 mask_rev_in[4] input30/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyb_1
Xinput63 mgmt_gpio_in[34] input63/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
Xinput41 mgmt_gpio_in[14] input41/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyb_1
Xinput52 mgmt_gpio_in[24] input52/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyb_1
X_4583_ _4454_/Z _4583_/A2 _4583_/B _7396_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
Xhold803 _7961_/Q hold803/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
X_7371_ _7371_/D _7875_/RN _7410_/CLK _7371_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
Xinput96 wb_adr_i[10] input96/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_115_222 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6322_ _4460_/Z _6332_/A2 _6322_/B _7792_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
Xinput85 spimemio_flash_io0_do input85/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyb_1
Xhold825 _7636_/Q hold825/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
Xhold814 _7473_/Q hold814/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
Xinput74 pad_flash_io1_di _3664_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyb_1
Xhold836 _7408_/Q hold836/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
XFILLER_116_767 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6253_ hold585/Z _6264_/A2 _6254_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
Xhold847 _7363_/Q hold847/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
Xhold858 _7404_/Q hold858/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
Xhold869 _7386_/Q hold869/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
XFILLER_170_394 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5204_ _5338_/A1 _5663_/A1 _5381_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_103_428 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6184_ _7728_/Q _6191_/A2 _6185_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_130_247 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5135_ _5643_/A2 _5783_/A2 _5765_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_5066_ _5254_/A2 _5448_/A1 _5066_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_123_27 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_84_389 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4017_ _7616_/Q _5937_/A1 _4219_/A2 input16/Z hold55/I _7379_/Q _4020_/A2 VDD VSS
+ gf180mcu_fd_sc_mcu7t5v0__aoi222_1
XFILLER_72_507 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_38_751 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_65_570 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_37_283 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_53_721 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_16_69 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_25_467 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5968_ _4481_/I _5970_/A2 _5968_/B _7626_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_4919_ _5199_/B _5369_/B _4919_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__and2_2
XFILLER_166_601 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7707_ _7707_/D _7923_/RN _7816_/CLK _7707_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_138_325 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5899_ hold293/Z _5902_/A2 hold294/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_165_144 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_120_6 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7638_ _7638_/D input75/Z _7638_/CLK _7638_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffsnq_1
XFILLER_107_712 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7569_ _7569_/D input75/Z _7638_/CLK _7569_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffsnq_1
XFILLER_134_531 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_134_575 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_88_662 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_88_673 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_102_494 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_28_250 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_16_412 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_43_286 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_12_673 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_12_662 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_157_667 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_144_328 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_156_188 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_125_564 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_140_534 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_415 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_404 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_112_258 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_112_247 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_448 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_437 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_426 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_459 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_121_792 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_93_131 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_94_676 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6940_ _6950_/A1 _6950_/A2 _6941_/A2 _7207_/B1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor3_4
XFILLER_54_507 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_81_337 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_19_283 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_47_570 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_19_294 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6871_ _6871_/A1 _6871_/A2 _6871_/A3 _6872_/C VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand3_1
X_5822_ hold646/Z _5827_/A2 _5823_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_35_798 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5753_ _5099_/B _5753_/A2 _5753_/B _5753_/C _5800_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_22_437 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_50_757 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_147_100 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4704_ _3819_/Z hold16/Z _4705_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_148_656 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_147_133 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_147_144 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5684_ _5701_/C _5684_/A2 _5684_/A3 _5684_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__and3_1
X_4635_ hold467/Z _3830_/Z _4635_/B hold468/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_7423_ _7423_/D _7901_/RN _7849_/CLK _7997_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_108_509 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_163_637 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
Xhold600 _7712_/Q hold600/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
Xhold611 _7794_/Q hold611/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
XFILLER_116_531 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7354_ _7354_/D _7961_/RN _7531_/CLK _7354_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffsnq_1
X_4566_ _6539_/A1 _4568_/A2 _4566_/B _7389_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
Xhold644 _7634_/Q hold644/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
Xmax_cap352 _5433_/C _5422_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__buf_4
XFILLER_118_49 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6305_ _4460_/Z _6315_/A2 _6305_/B _7784_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
Xhold622 hold622/I _7684_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
Xhold633 hold633/I _7365_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
Xhold688 _7808_/Q hold688/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
Xhold655 hold655/I _6096_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
Xhold677 _7880_/Q hold677/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
X_4497_ hold517/Z _4504_/A2 hold518/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_7285_ _7285_/A1 _7285_/A2 _7289_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
Xhold666 _7700_/Q hold666/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
X_6236_ hold16/Z hold6/Z _6236_/B hold58/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_131_567 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xhold699 _7649_/Q hold699/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
XFILLER_134_37 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6167_ hold524/Z _6174_/A2 _6168_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_69_150 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_960 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_971 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_5118_ _5309_/A1 _3723_/I _4898_/Z _5689_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand3_4
XFILLER_94_19 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_84_120 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_982 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_993 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_57_323 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_57_334 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6098_ hold64/Z _6106_/A2 _6098_/B hold112/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_84_131 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_73_805 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_5049_ _5309_/A1 _3723_/I _5006_/B _5448_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor3_4
XFILLER_26_732 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_27_79 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_26_798 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_43_23 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_80_392 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_13_459 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_25_286 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_43_34 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_21_481 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_40_289 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_111_2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_162_681 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_4_179 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_4_17 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_122_534 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_68_64 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_352 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_363 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_76_632 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_48_312 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_91_602 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_84_41 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_76_687 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_76_676 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_48_356 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_48_367 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_29_570 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_48_389 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_84_96 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_63_348 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_16_264 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_17_798 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_177_707 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_71_392 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_270 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_292 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_281 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_129_111 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_129_122 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_83_6 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_12_481 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_31_278 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_129_144 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_8_463 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_69_4 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4420_ _4420_/I _4420_/ZN VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_160_629 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4351_ _4331_/Z _6622_/A2 _6569_/A3 _4361_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor3_2
XFILLER_113_545 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_113_534 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_99_779 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7070_ _7882_/Q _7203_/B1 _7204_/A2 _7842_/Q _7834_/Q _7203_/A2 _7077_/A1 VDD VSS
+ gf180mcu_fd_sc_mcu7t5v0__aoi222_1
X_4282_ _4282_/A1 _4282_/A2 _4283_/A4 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_113_567 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_98_267 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_86_429 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_86_418 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_86_407 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6021_ _6553_/A1 _6021_/A2 _6021_/B hold120/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_104_29 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_82_602 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_39_345 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7972_ _7972_/D _7325_/Z _7972_/CLK hold1/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_94_495 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_82_624 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6923_ _7914_/Q _7913_/Q _6950_/A1 _6955_/A4 _7201_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor4_4
XFILLER_70_808 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_66_197 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_62_392 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6854_ _7401_/Q _6893_/A2 _6890_/B1 _7395_/Q _6867_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_167_228 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5805_ _5805_/A1 _5804_/Z _5805_/B _5806_/A4 VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_6785_ _7721_/Q _6881_/A2 _6882_/B1 _7657_/Q _6787_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_3997_ _7883_/Q _6503_/A1 _4232_/A2 input8/Z _3997_/C _3998_/A4 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi221_1
XFILLER_23_779 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5736_ _5736_/A1 _5736_/A2 _5706_/Z _5736_/A4 _5785_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand4_1
XFILLER_182_209 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5667_ _5667_/A1 _5602_/Z _5667_/A3 _5748_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_175_283 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_148_486 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_89_19 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4618_ _4454_/Z _4618_/A2 _4618_/B _7410_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_7406_ _7406_/D _7875_/RN _7822_/CLK _7406_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
X_5598_ _5087_/C _5579_/B _5777_/A2 _5777_/A1 _5665_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_7337_ _7337_/D _7292_/Z _4415_/A2 _7337_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_150_128 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
Xhold463 hold463/I _7825_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
XFILLER_89_212 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xhold430 _7640_/Q hold430/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
Xhold441 _7882_/Q hold441/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
Xhold452 _8002_/I hold452/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
X_4549_ _4549_/A1 _6537_/A2 _4553_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_7268_ _7268_/A1 _7277_/B _7268_/B _7955_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_150_139 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_145_69 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
Xhold496 hold496/I _7708_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
Xhold485 hold485/I _7420_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
XFILLER_104_534 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
Xhold474 hold474/I _4519_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
X_6219_ hold16/Z _6225_/A2 _6219_/B hold44/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_38_34 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7199_ _7199_/A1 _7199_/A2 _7198_/Z _7209_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_85_451 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_38_67 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_790 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_58_676 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_173_4 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1901 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_73_668 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_72_134 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_45_337 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_45_348 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1934 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1923 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1912 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_60_318 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_159_707 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_159_2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1967 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1956 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1945 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_13_212 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1989 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1978 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_41_565 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_167_773 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_166_250 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_127_637 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_182_754 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_181_286 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_123_810 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_5_499 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_5_488 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_135_692 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_150_662 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_95_215 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_135_80 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_95_73 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_64_602 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_193 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_48_120 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_91_410 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_64_624 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_17_540 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3920_ _7976_/Q _7413_/Q _4427_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_4
XFILLER_17_551 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_51_318 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_44_392 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3851_ hold76/Z hold82/Z _6350_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_4
X_3782_ hold49/I hold24/Z hold25/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_20_727 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_20_738 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6570_ _7905_/Q _6570_/A2 _6570_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_5521_ _5521_/A1 _5521_/A2 _5522_/B2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_118_615 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_74_2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_9_761 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_157_283 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_157_294 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_9_783 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_8_260 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_145_456 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5452_ _4993_/C _5527_/A1 _5543_/C _5452_/C _5454_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XFILLER_117_136 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_173_798 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_5383_ _5576_/B2 _5382_/Z _5565_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_132_117 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_4403_ _7334_/Q input38/Z _4403_/B _7979_/Q _4404_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi211_1
X_4334_ _7630_/Q _4335_/A2 _4334_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__and2_4
X_7122_ _7828_/Q _7202_/A2 _7202_/B1 _7788_/Q _7764_/Q _7202_/C2 _7129_/A1 VDD VSS
+ gf180mcu_fd_sc_mcu7t5v0__aoi222_1
XFILLER_115_17 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_7053_ _7053_/A1 _7053_/A2 _7053_/A3 _7053_/A4 _7054_/A4 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand4_1
XFILLER_140_161 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6004_ _6553_/A1 _6004_/A2 _6004_/B hold209/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_86_237 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_4265_ _7569_/Q _5841_/A1 _4599_/A1 _7403_/Q _4267_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_4196_ _7557_/Q _5812_/A1 _4754_/A1 _7467_/Q _4198_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_82_454 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_7955_ _7955_/D _7959_/RN _4411_/I1 _7955_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XTAP_1219 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1208 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_70_605 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_42_318 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6906_ _6599_/Z _6950_/A2 _6941_/A2 _7189_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor3_4
XFILLER_70_638 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7886_ _7886_/D _7900_/RN _7900_/CLK _7886_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffsnq_1
XFILLER_168_504 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6837_ _7723_/Q _6881_/A2 _6881_/B1 _7699_/Q _6839_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_148_250 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6768_ _7624_/Q _6659_/Z _6884_/B1 _7688_/Q _6771_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_164_732 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5719_ _5719_/A1 _5677_/Z _5719_/A3 _5719_/A4 _7542_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__or4_1
XFILLER_108_114 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6699_ _7645_/Q _6880_/C2 _6881_/B1 _7693_/Q _7807_/Q _6880_/B1 _6702_/A1 VDD VSS
+ gf180mcu_fd_sc_mcu7t5v0__aoi222_1
XFILLER_136_445 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_164_798 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_163_286 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_108_169 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
Xhold271 _7457_/Q hold271/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
XFILLER_117_692 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
Xhold260 _7829_/Q hold260/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
XFILLER_132_673 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xhold293 _8004_/I hold293/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
XFILLER_78_705 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
Xhold282 hold282/I _7884_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
XFILLER_2_458 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_49_33 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_172_34 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_77_215 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_58_440 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_65_32 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_46_602 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_46_635 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_18_348 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1742 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1731 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1720 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_61_638 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_26_392 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1775 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1764 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1753 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_14_543 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1797 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1786 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_167_570 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_139_283 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_182_562 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_6_742 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_155_798 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_5_241 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_107_180 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_46_6 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4050_ _7873_/Q _6486_/A1 _6039_/A1 hold79/I _6022_/A1 _7655_/Q _4052_/A2 VDD VSS
+ gf180mcu_fd_sc_mcu7t5v0__aoi222_1
XFILLER_49_451 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_110_389 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xinput6 mask_rev_in[11] input6/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XFILLER_49_462 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_37_679 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_52_605 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4952_ _5496_/A1 _5741_/A1 _5602_/A1 _7518_/Q _5474_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai31_1
X_7740_ _7740_/D _7877_/RN _7773_/CLK _7740_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffsnq_1
XFILLER_51_104 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3903_ _7877_/Q _6486_/A1 _6005_/A1 _7651_/Q _6520_/A1 _7893_/Q _3906_/A2 VDD VSS
+ gf180mcu_fd_sc_mcu7t5v0__aoi222_1
X_7671_ _7671_/D _7923_/RN _7735_/CLK _7671_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
X_4883_ _4883_/A1 _7285_/A2 _4887_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_3834_ hold609/Z hold89/Z _5886_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_4
X_6622_ _6622_/A1 _6622_/A2 _6622_/B _7919_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_3765_ _3765_/A1 _3765_/A2 _3765_/B _7973_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_6553_ _6553_/A1 _6553_/A2 _6553_/B hold270/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_173_540 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_173_551 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5504_ _5545_/A2 _5687_/B _5504_/A3 _5504_/B1 _5543_/B _5505_/A4 VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai32_1
XFILLER_146_743 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_118_456 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3696_ _7735_/Q _3696_/ZN VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_6484_ hold239/Z _6485_/A2 hold240/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_145_286 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5435_ _5435_/A1 _5435_/A2 _5446_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_10_27 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
Xoutput310 _7941_/Q wb_ack_o VDD VSS gf180mcu_fd_sc_mcu7t5v0__buf_4
XFILLER_160_212 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xoutput332 _7947_/Q wb_dat_o[29] VDD VSS gf180mcu_fd_sc_mcu7t5v0__buf_4
Xoutput321 _7481_/Q wb_dat_o[19] VDD VSS gf180mcu_fd_sc_mcu7t5v0__buf_4
X_5366_ _4965_/B _5366_/A2 _4993_/C _5689_/A1 _5622_/A1 _5572_/C VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai32_1
X_4317_ _7414_/Q _4294_/Z _4317_/A3 _4318_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor3_1
X_5297_ _5006_/C _5709_/A2 _5297_/B _5378_/C _5299_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi211_1
X_7105_ _7105_/A1 _7105_/A2 _7105_/A3 _7105_/A4 _7106_/A4 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand4_1
XFILLER_59_215 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7036_ _7849_/Q _7193_/A2 _7189_/A2 hold84/I _7203_/B1 _7881_/Q _7039_/A2 VDD VSS
+ gf180mcu_fd_sc_mcu7t5v0__aoi222_1
XFILLER_68_760 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4248_ _4248_/A1 _4248_/A2 _4248_/A3 _4248_/A4 _4283_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand4_2
XFILLER_142_37 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_28_602 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_55_410 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_16_808 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4179_ _4179_/A1 _4179_/A2 _4179_/A3 _4179_/A4 _4187_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand4_1
XFILLER_35_24 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_7938_ _7938_/D _7938_/RN _7938_/CLK _7938_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_15_329 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_42_126 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_43_638 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1005 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1016 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1038 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1027 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1049 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_7869_ _7869_/D _7901_/RN _7869_/CLK _7869_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_168_389 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_149_570 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_164_540 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_137_798 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_3_712 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_151_212 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_124_448 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_4_2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_120_621 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_116_71 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_120_676 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_76_64 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_65_207 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_59_760 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_46_410 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_46_421 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_58_281 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_74_763 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_34_605 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2262 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2251 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2240 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_61_424 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2295 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2284 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2273 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
Xclkbuf_leaf_41_csclk clkbuf_3_7__f_csclk/Z _7747_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XTAP_1550 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1594 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1583 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1572 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1561 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_660 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_90 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_159_367 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_41_192 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_42_693 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
Xclkbuf_leaf_56_csclk clkbuf_3_6__f_csclk/Z _7792_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_155_540 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_155_595 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5220_ _5538_/A1 _5042_/Z _5176_/B _5652_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_127_286 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_115_437 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5151_ _5151_/A1 _5151_/A2 _5024_/Z _5539_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_142_278 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_96_321 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_37_2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5082_ _5319_/C _5714_/B1 _5307_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_4102_ _7808_/Q _6350_/A1 _4232_/A2 input5/Z _6418_/A1 _7840_/Q _4104_/A3 VDD VSS
+ gf180mcu_fd_sc_mcu7t5v0__aoi222_1
X_4033_ _7664_/Q _6039_/A1 _4505_/A1 _7367_/Q _6333_/A1 _7802_/Q _4035_/A3 VDD VSS
+ gf180mcu_fd_sc_mcu7t5v0__aoi222_1
XFILLER_49_281 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_80_744 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_25_638 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5984_ hold644/Z _5987_/A2 _5985_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_7723_ _7723_/D _7853_/RN _7811_/CLK _7723_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
X_4935_ _5230_/A1 _5271_/A3 _5482_/B2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_2
XFILLER_80_788 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_21_811 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_33_682 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_178_676 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7654_ _7654_/D _7923_/RN _7734_/CLK _7654_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffsnq_1
XFILLER_20_321 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4866_ hold891/Z _4867_/A2 hold892/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_138_529 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3817_ hold27/Z _4686_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_7585_ _7585_/D _7923_/RN _7698_/CLK _7585_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
X_6605_ _7914_/Q _7913_/Q _6950_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_4
X_4797_ _7230_/A1 _4795_/S _4797_/B _7485_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_181_808 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3748_ _7344_/Q _7411_/Q _3751_/A2 _3749_/S VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_119_765 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_6536_ _6553_/A1 _6536_/A2 _6536_/B hold257/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_180_318 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_119_798 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_133_212 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6467_ hold242/Z _6468_/A2 hold243/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_97_19 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3679_ hold98/I _3679_/ZN VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_5418_ _5692_/B _5563_/B2 _5618_/A3 _5419_/C VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor3_1
X_6398_ hold233/Z _6400_/A2 _6398_/B hold290/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
Xoutput195 _3681_/ZN mgmt_gpio_oeb[31] VDD VSS gf180mcu_fd_sc_mcu7t5v0__buf_4
XFILLER_153_25 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5349_ _5482_/B2 _5510_/A2 _5493_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
Xoutput173 _3701_/ZN mgmt_gpio_oeb[11] VDD VSS gf180mcu_fd_sc_mcu7t5v0__buf_4
Xoutput184 _3691_/ZN mgmt_gpio_oeb[21] VDD VSS gf180mcu_fd_sc_mcu7t5v0__buf_4
XFILLER_0_737 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_87_354 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_102_687 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_102_676 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7019_ _7880_/Q _7203_/B1 _7204_/A2 _7840_/Q _7832_/Q _7203_/A2 _7025_/A1 VDD VSS
+ gf180mcu_fd_sc_mcu7t5v0__aoi222_1
XFILLER_46_34 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_16_605 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_28_498 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_70_254 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_102_84 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_62_33 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_12_811 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_141_2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_11_343 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_109_231 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_11_398 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_171_307 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_164_392 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_125_757 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_109_286 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_11_70 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_127_92 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_608 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_619 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_78_321 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_93_302 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_93_357 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_34_402 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2070 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2092 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2081 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_62_788 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_1391 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1380 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_4720_ hold767/Z _4731_/A2 _4721_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_174_112 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4651_ hold271/Z _3830_/Z _4651_/B _4652_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_147_348 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_128_540 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
Xinput20 mask_rev_in[24] input20/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyb_1
Xinput31 mask_rev_in[5] input31/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyb_1
Xinput64 mgmt_gpio_in[35] input64/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XFILLER_162_318 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xinput42 mgmt_gpio_in[15] input42/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyb_1
Xinput53 mgmt_gpio_in[25] input53/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyb_1
X_7370_ _7370_/D input75/Z _7875_/CLK _7370_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffsnq_1
X_4582_ hold839/Z _4583_/A2 _4583_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
Xinput97 wb_adr_i[11] input97/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_115_212 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6321_ hold645/Z _6332_/A2 _6322_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
Xinput86 spimemio_flash_io0_oeb input86/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyb_1
Xhold826 _7999_/I hold826/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
Xhold837 _7505_/Q hold837/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
XFILLER_6_380 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xinput75 porb input75/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__buf_16
Xhold815 _7757_/Q hold815/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
Xhold804 _7895_/Q hold804/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
XFILLER_170_340 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
Xhold848 hold848/I _4507_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
Xhold859 _7410_/Q hold859/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
X_6252_ _4454_/Z _6264_/A2 _6252_/B _7759_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_5203_ _5203_/I _5375_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_6183_ hold64/Z _6191_/A2 _6183_/B _7727_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_5134_ _3723_/I _5777_/A1 _5538_/A1 _5026_/Z _5451_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__and4_1
XFILLER_97_641 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_69_354 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5065_ _5476_/B _5689_/A1 _5072_/B _5359_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_111_495 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_96_195 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_4016_ _4013_/Z _4016_/A2 _4016_/A3 _4025_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_16_37 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_80_585 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5967_ hold658/Z _5970_/A2 _5968_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_4918_ _3722_/I _5006_/B _5006_/C _3728_/I _4945_/B1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand4_1
X_7706_ _7706_/D _7938_/RN _7738_/CLK _7706_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
X_5898_ _6549_/A1 _5902_/A2 _5898_/B _7593_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_21_641 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7637_ _7637_/D input75/Z _7637_/CLK _7637_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffsnq_1
XFILLER_166_657 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_166_646 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_119_540 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4849_ hold408/Z _4852_/A2 _4850_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_119_551 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_7568_ _7568_/D _7875_/RN _7874_/CLK _7568_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_181_638 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_146_392 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_134_510 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_113_6 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6519_ _6553_/A1 _6519_/A2 _6519_/B hold267/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_7499_ _7499_/D _7503_/CLK _7499_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_107_779 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_106_256 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_134_598 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_122_727 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_121_215 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_589 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_180_34 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_48_538 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_75_357 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_28_240 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_90_338 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_73_32 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_44_744 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_44_766 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_71_574 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_157_635 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_129_304 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_172_605 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_11_195 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_7_144 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_171_137 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_125_554 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_98_51 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_180_693 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_405 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_79_641 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_449 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_438 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_427 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_416 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_93_121 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_82_806 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_54_519 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_93_176 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_35_722 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_62_530 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6870_ _7960_/Q _6880_/A2 _6893_/C1 _7472_/Q _6871_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_179_215 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_62_563 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5821_ _4454_/Z _5827_/A2 _5821_/B _7559_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_5752_ _5777_/A1 _5608_/B _5752_/B1 _4996_/Z _5752_/C _5753_/C VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi221_1
XFILLER_15_490 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_50_747 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_148_602 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4703_ hold320/Z _4718_/A1 hold321/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_148_646 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5683_ _5433_/C _5683_/A2 _5684_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_30_460 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_163_616 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4634_ _3830_/Z hold64/I _4635_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_7422_ _7422_/D _7901_/RN _7422_/CLK _7996_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
Xhold612 _7986_/I hold612/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
Xhold601 hold601/I _6151_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
XFILLER_118_17 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7353_ _7353_/D _7961_/RN _7531_/CLK _7353_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffsnq_1
X_4565_ hold753/Z _4568_/A2 _4566_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_128_392 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
Xmax_cap353 _7877_/RN _7853_/RN VDD VSS gf180mcu_fd_sc_mcu7t5v0__buf_20
Xhold645 _7792_/Q hold645/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
Xhold634 _7678_/Q hold634/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
X_6304_ hold685/Z _6315_/A2 _6305_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
Xhold623 _7357_/Q hold623/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
X_7284_ _7284_/I _7959_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_171_682 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
Xhold678 _7662_/Q hold678/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
XFILLER_103_215 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
Xhold656 hold656/I _7686_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
X_4496_ _6545_/A1 _4504_/A2 _4496_/B hold249/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
Xhold667 hold667/I _6126_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
Xhold689 _7377_/Q hold689/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
X_6235_ hold57/Z hold6/Z _6236_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_6166_ hold64/Z _6174_/A2 _6166_/B hold91/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_97_460 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_950 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_961 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_5117_ _5392_/A1 _5344_/A2 _5680_/B2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_2
X_6097_ hold110/Z _6106_/A2 hold111/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_972 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_983 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_994 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_5048_ _5309_/A1 _3723_/I _5254_/A2 _5102_/B1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor3_1
XFILLER_111_292 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_57_357 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_150_37 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_26_744 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_40_202 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_53_585 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6999_ _7775_/Q _7200_/A2 _7201_/A2 _7749_/Q _7200_/B1 _7863_/Q _7000_/A4 VDD VSS
+ gf180mcu_fd_sc_mcu7t5v0__aoi222_1
XFILLER_159_57 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_138_101 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_178_281 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_139_635 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_154_616 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_154_605 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_126_318 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_21_493 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_175_34 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_5_637 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_104_2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_162_693 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_162_671 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_107_576 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_68_43 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_68_54 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_48_302 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_49_803 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_124_60 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_75_154 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_84_53 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_75_165 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_90_179 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_17_766 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_140_92 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_32_736 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_32_747 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_260 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_129_101 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_293 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_282 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_271 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_129_134 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_12_460 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_8_453 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_4350_ _6567_/A1 _7905_/Q _6569_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_141_800 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_140_321 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_125_384 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_113_557 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4281_ _4281_/A1 _4281_/A2 _4281_/A3 _4281_/A4 _4282_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor4_1
XFILLER_101_708 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6020_ hold119/Z _6021_/A2 _6021_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_79_493 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_94_463 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_39_357 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_55_806 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_7971_ _7971_/D _7324_/Z _7972_/CLK _7971_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_66_176 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xclkbuf_3_3__f_csclk clkbuf_0_csclk/Z clkbuf_3_3__f_csclk/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_54_305 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_54_316 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6922_ _6599_/Z _6955_/A4 _6908_/Z _7191_/B1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor3_4
XFILLER_120_29 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6853_ _7533_/Q _6878_/A2 _6853_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__or2_1
XFILLER_35_574 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5804_ _5804_/A1 _5804_/A2 _5804_/A3 _5804_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__or3_1
X_6784_ _7649_/Q _6880_/C2 _6882_/A2 _7380_/Q _7819_/Q _6880_/A2 _6787_/A1 VDD VSS
+ gf180mcu_fd_sc_mcu7t5v0__aoi222_1
X_3996_ _3996_/A1 _3996_/A2 _3996_/A3 _3997_/C VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_10_408 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5735_ _5104_/B _5735_/A2 _5247_/B _5724_/B _5735_/C _5736_/A4 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi221_1
XFILLER_31_780 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_136_605 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5666_ _5666_/A1 _5709_/A1 _5777_/A2 _5667_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_109_808 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_175_295 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_129_690 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_108_318 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4617_ hold859/Z _4618_/A2 _4618_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_7405_ _7405_/D _7875_/RN _7822_/CLK _7405_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
Xhold420 _7454_/Q hold420/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
X_5597_ _5417_/I _5450_/C _5656_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_7336_ _7336_/D _7291_/Z _4415_/A2 _7336_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_144_671 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4548_ _6553_/A1 _4548_/A2 _4548_/B _7382_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
Xhold431 hold431/I _5998_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
Xhold442 hold442/I _6513_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
Xhold453 hold453/I _5896_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
X_7267_ _7267_/A1 _7280_/A2 _7277_/B _7267_/C _7268_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi211_1
Xhold464 _7461_/Q hold464/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
X_4479_ hold49/Z _7273_/A1 _4480_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
Xhold486 _7748_/Q hold486/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
Xhold475 hold475/I _7369_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
X_6218_ _7744_/Q _6225_/A2 _6219_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_131_354 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xhold497 _7706_/Q hold497/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
X_7198_ _7198_/A1 _7198_/A2 _7198_/A3 _7198_/A4 _7198_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__and4_1
XFILLER_58_611 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_58_622 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6149_ hold64/Z _6157_/A2 hold85/Z hold86/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
XTAP_780 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_791 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_161_69 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_85_496 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1924 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1913 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1902 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_72_179 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_54_34 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1968 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1957 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1946 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1935 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_14_747 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1979 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_70_44 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_70_33 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_9_239 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_167_763 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_119_82 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_181_298 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_122_321 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_96_717 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_135_70 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_95_30 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_89_780 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_76_452 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_76_441 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_49_666 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_76_463 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_48_176 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_48_187 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_51_308 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_91_499 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3850_ hold53/Z _3864_/A2 hold81/Z _3864_/A4 hold82/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand4_4
X_3781_ hold192/Z hold87/Z _7414_/Q _3781_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_20_717 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_32_577 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_32_588 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_32_599 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5520_ _5359_/B _5520_/A2 _5520_/B _5520_/C _5522_/B1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XFILLER_118_605 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_172_210 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_117_115 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_8_250 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_173_777 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5451_ _5774_/A1 _5643_/A2 _5451_/B _5460_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_67_2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5382_ _5022_/B _5205_/Z _5382_/A3 _5382_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__or3_1
X_4402_ _4402_/A1 _4334_/Z _4402_/B _7334_/Q _4403_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XFILLER_99_511 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_153_490 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_141_641 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_113_310 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_99_522 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4333_ input67/Z _7582_/Q _4335_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_2
X_7121_ _7121_/A1 _7121_/A2 _7121_/A3 _7121_/A4 _7130_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand4_1
XFILLER_113_354 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_101_505 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7052_ hold78/I _7195_/A2 _7190_/B1 _7615_/Q _7053_/A4 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_5_83 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4264_ _4264_/A1 _4264_/A2 _4264_/A3 _4264_/A4 _4281_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand4_1
X_6003_ hold207/Z _6004_/A2 hold208/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_39_132 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4195_ _7775_/Q _6282_/A1 _4888_/A1 _7536_/Q _6401_/A1 _7831_/Q _4198_/A2 VDD VSS
+ gf180mcu_fd_sc_mcu7t5v0__aoi222_1
XFILLER_95_783 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7954_ _7954_/D _7959_/RN _7959_/CLK _7954_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_82_444 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_27_327 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_43_809 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6905_ _6905_/A1 _6905_/A2 _6941_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_4
XTAP_1209 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_54_179 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_7885_ _7885_/D _7901_/RN _7901_/CLK _7885_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_24_15 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6836_ _7821_/Q _6880_/A2 _6880_/B1 _7813_/Q _7651_/Q _6880_/C2 _6839_/A1 VDD VSS
+ gf180mcu_fd_sc_mcu7t5v0__aoi222_1
XFILLER_24_37 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_6767_ _7736_/Q _6830_/B _6889_/A2 _7704_/Q _6767_/C _6771_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi221_1
XFILLER_10_205 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5718_ _5590_/B _5581_/B _5718_/A3 _5719_/A4 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor3_1
X_3979_ _7811_/Q _6350_/A1 _6333_/A1 _7803_/Q _3992_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_164_722 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_148_262 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_109_638 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6698_ _7637_/Q _6890_/A2 _6665_/Z _7741_/Q _6698_/C _6707_/B1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi221_1
XFILLER_164_744 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5649_ _5673_/A3 _5647_/B _5649_/A3 _5649_/A4 _5655_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand4_1
XFILLER_108_148 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_108_126 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_40_69 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_123_118 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7319_ _7877_/RN _4334_/Z _7319_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_123_129 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_117_682 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
Xhold261 hold261/I _6400_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
XFILLER_104_321 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
Xhold250 _7845_/Q hold250/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
Xhold272 _4741_/Z _7457_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
Xhold294 hold294/I _5900_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
Xhold283 _7844_/Q hold283/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
XFILLER_93_709 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_19_806 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_105_73 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_58_463 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_58_485 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2400 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_171_2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1743 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1732 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1721 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1710 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_73_499 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_60_105 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1776 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1765 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1754 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1798 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1787 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_14_599 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_41_352 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_127_424 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_154_254 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_170_747 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_5_286 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_123_641 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_150_460 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_83_208 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_77_783 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xinput7 mask_rev_in[12] input7/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XFILLER_37_614 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_92_742 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_92_731 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_76_271 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_64_433 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_49_496 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4951_ _4951_/A1 _4951_/A2 _4951_/B _5016_/B _5602_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai211_4
XFILLER_36_179 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_3902_ _7885_/Q _6503_/A1 _5903_/A1 input42/Z _4231_/B1 input70/Z _3906_/A1 VDD VSS
+ gf180mcu_fd_sc_mcu7t5v0__aoi222_1
X_7670_ _7670_/D _7923_/RN _7734_/CLK _7670_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffsnq_1
X_4882_ _4454_/Z _4882_/A2 _4882_/B hold821/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_3833_ _3783_/Z _3925_/A2 hold75/Z _3963_/A4 hold89/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand4_4
X_6621_ _7919_/Q _6621_/A2 _6622_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_177_379 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_177_357 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3764_ _3765_/A2 _3764_/A2 _3765_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_6552_ hold268/Z _6553_/A2 hold269/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_9_570 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3695_ hold68/I _3695_/ZN VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_5503_ _5797_/A2 _5546_/A2 _5546_/B1 _5543_/B _5503_/C _5509_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai221_1
X_6483_ hold233/Z _6485_/A2 _6483_/B hold301/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_5434_ _5789_/A1 _5614_/A3 _5625_/A2 _5434_/A4 _5435_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand4_1
Xoutput300 _4331_/Z serial_clock VDD VSS gf180mcu_fd_sc_mcu7t5v0__buf_4
XFILLER_114_630 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
Xoutput322 _7497_/Q wb_dat_o[1] VDD VSS gf180mcu_fd_sc_mcu7t5v0__buf_4
Xoutput333 _7498_/Q wb_dat_o[2] VDD VSS gf180mcu_fd_sc_mcu7t5v0__buf_4
Xoutput311 _7496_/Q wb_dat_o[0] VDD VSS gf180mcu_fd_sc_mcu7t5v0__buf_4
XFILLER_160_268 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5365_ _5797_/A1 _5099_/B _5365_/B1 _5681_/A1 _5408_/C VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai22_1
X_7104_ _7883_/Q _7203_/B1 _7204_/A2 _7843_/Q _7105_/A4 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_4316_ _7337_/Q _7336_/Q hold87/I _4317_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_5296_ _5371_/C _5405_/B _5378_/C VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_141_471 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7035_ _7035_/A1 _7035_/A2 _7035_/A3 _7035_/A4 _7035_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__and4_1
XFILLER_101_357 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_101_346 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_75_709 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4247_ _7676_/Q _6073_/A1 _5971_/A1 _7628_/Q _4248_/A4 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_142_27 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4178_ _7759_/Q _6248_/A1 _4549_/A1 _7384_/Q _4179_/A4 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_83_753 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_82_252 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_27_168 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_55_477 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_7937_ _7937_/D _7938_/RN _7938_/CLK _7937_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XTAP_1028 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_105 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_42_116 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_55_499 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_1006 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1017 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_7868_ _7868_/D _7900_/RN _7878_/CLK _7868_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XTAP_1039 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_6819_ _6819_/A1 _6819_/A2 _6819_/A3 _6819_/A4 _6825_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand4_1
XFILLER_23_352 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_51_672 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7799_ _7799_/D _7875_/RN _7863_/CLK _7799_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffsnq_1
XFILLER_51_35 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_109_424 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_137_766 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_109_479 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_152_747 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_152_769 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_105_641 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_3_779 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_132_460 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_104_151 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_116_83 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_76_32 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_59_783 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_74_742 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_18_124 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_73_241 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2252 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2241 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2230 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_92_53 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_73_296 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_18_179 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2296 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2285 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2274 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2263 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1551 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1540 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_14_330 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1584 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1573 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1562 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_30_812 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_80 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_91 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_159_357 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_147_508 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_1595 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_174_327 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_128_744 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_155_563 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_157_90 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_127_298 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5150_ _5151_/A1 _5151_/A2 _5024_/Z _5150_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__and3_1
XFILLER_151_780 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_97_812 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5081_ _4898_/Z _5254_/A3 _5714_/B1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_2
X_4101_ input37/Z _5903_/A1 _4488_/A1 _7357_/Q _5874_/A1 _7583_/Q _4104_/A2 VDD VSS
+ gf180mcu_fd_sc_mcu7t5v0__aoi222_1
XFILLER_57_709 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4032_ _4032_/A1 _4032_/A2 _4036_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_37_400 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_110_176 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_92_561 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_92_550 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_65_753 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_5983_ _4476_/I _5987_/A2 _5983_/B _7633_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_18_680 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_24_105 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_37_499 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_178_600 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7722_ _7722_/D _7853_/RN _7722_/CLK _7722_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
X_4934_ _5199_/B _5201_/B _5271_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_4
X_4865_ hold47/Z _4867_/A2 _4865_/B hold404/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_20_311 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_7653_ _7653_/D _7938_/RN _7653_/CLK _7653_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffsnq_1
XFILLER_177_176 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3816_ hold26/Z _3925_/A2 hold75/I hold71/I hold27/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__or4_4
X_7584_ _7584_/D _7923_/RN _7698_/CLK _7584_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
X_6604_ _7913_/Q _6609_/A2 _6604_/B _7913_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_4796_ _7485_/Q _4795_/S _4797_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_3747_ _4284_/A1 _3763_/B _3747_/B _7977_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_118_210 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6535_ hold255/Z _6536_/A2 hold256/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_3678_ _7873_/Q _3678_/ZN VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_146_596 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_134_747 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_133_224 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_106_427 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6466_ hold233/Z _6468_/A2 _6466_/B hold298/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_5417_ _5417_/I _5446_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_6397_ hold288/Z _6400_/A2 hold289/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
Xoutput174 _3700_/ZN mgmt_gpio_oeb[12] VDD VSS gf180mcu_fd_sc_mcu7t5v0__buf_4
XFILLER_114_460 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xoutput185 _3690_/ZN mgmt_gpio_oeb[22] VDD VSS gf180mcu_fd_sc_mcu7t5v0__buf_4
XFILLER_102_611 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5348_ _5685_/B _5624_/A2 _5642_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_88_812 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_87_311 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xoutput196 _3680_/ZN mgmt_gpio_oeb[32] VDD VSS gf180mcu_fd_sc_mcu7t5v0__buf_4
X_7018_ _7750_/Q _7201_/A2 _7201_/B1 _7670_/Q _7023_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_5279_ _5616_/A1 _5237_/Z _5712_/B _5573_/B _5282_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XFILLER_75_539 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_68_591 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_46_24 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_71_723 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_71_734 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_71_712 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_102_52 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_31_609 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_169_633 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_169_611 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_70_277 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_30_108 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_178_34 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_168_176 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_134_2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_156_338 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_140_717 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_112_419 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_97_119 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_97_108 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_79_812 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_609 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_87_64 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_39_709 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_120_463 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_59_591 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_59_580 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_81_509 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_19_455 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_19_499 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2060 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2093 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2082 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2071 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1392 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1381 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1370 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_159_176 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4650_ _3830_/Z hold2/Z _4651_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_1
Xinput21 mask_rev_in[25] input21/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyb_1
Xinput10 mask_rev_in[15] input10/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XFILLER_174_179 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xinput43 mgmt_gpio_in[16] input43/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyb_1
Xinput54 mgmt_gpio_in[26] input54/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyb_1
Xinput32 mask_rev_in[6] input32/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyb_1
X_4581_ _6539_/A1 _4583_/A2 _4581_/B _7395_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_6320_ _4454_/Z _6332_/A2 _6320_/B _7791_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
Xinput65 mgmt_gpio_in[36] _8008_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyc_1
Xinput98 wb_adr_i[12] input98/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
Xhold827 _7709_/Q hold827/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
XFILLER_116_747 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
Xinput87 spimemio_flash_io1_do _8007_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyb_1
Xhold805 _7878_/Q hold805/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
Xinput76 qspi_enabled _4387_/S VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
Xhold816 _7384_/Q hold816/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
XFILLER_170_330 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_115_246 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_107_19 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_6_392 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xhold849 hold849/I _7363_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
Xhold838 _7400_/Q hold838/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
X_6251_ hold878/Z _6264_/A2 _6252_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_5202_ _5202_/A1 _5202_/A2 _5371_/B _5371_/C _5203_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_2
X_6182_ hold69/Z _6191_/A2 _6183_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_88_108 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5133_ _5309_/A1 _3723_/I _5394_/A1 _5006_/C _5645_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand4_4
XFILLER_123_290 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_69_333 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5064_ _5301_/A1 _5062_/Z _5064_/B _5072_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_97_697 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_84_336 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_84_325 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_29_219 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_57_528 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_57_539 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_84_347 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4015_ _7672_/Q _6056_/A1 _5886_/A1 input56/Z _5817_/A1 _7562_/Q _4016_/A3 VDD VSS
+ gf180mcu_fd_sc_mcu7t5v0__aoi222_1
XFILLER_25_425 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_53_712 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_80_531 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_12_108 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_5966_ _6549_/A1 _5970_/A2 _5966_/B _7625_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_25_469 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_52_266 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_53_789 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_4917_ _3722_/I _5006_/B _5006_/C _3728_/I _4917_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__and4_2
XFILLER_178_452 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7705_ _7705_/D _7923_/RN _7735_/CLK _7705_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
X_5897_ hold697/Z _5902_/A2 _5898_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_178_463 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7636_ _7636_/D input75/Z _7638_/CLK _7636_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffsnq_1
XFILLER_32_37 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_4848_ _4848_/A1 _6537_/A2 _4852_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_148_37 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_180_105 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7567_ _7567_/D _7875_/RN _7567_/CLK _7567_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffsnq_1
XFILLER_5_808 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4779_ _4779_/A1 _6537_/A2 _4783_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_107_725 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_6518_ hold265/Z _6519_/A2 hold266/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_4_318 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7498_ _7498_/D _7503_/CLK _7498_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_6449_ hold233/Z _6451_/A2 _6449_/B _7852_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_106_6 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xclkbuf_leaf_40_csclk clkbuf_3_7__f_csclk/Z _7809_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_122_717 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_115_780 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_88_620 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_524 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_102_463 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_88_686 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_87_163 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_87_141 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_579 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_57_34 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_102_496 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xclkbuf_leaf_55_csclk clkbuf_3_6__f_csclk/Z _7734_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_29_764 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_113_73 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_90_328 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_71_542 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_16_458 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_43_211 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_44_756 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_73_77 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_16_469 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_73_99 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_31_428 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_169_485 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_157_625 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_12_664 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_11_141 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_8_602 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_8_646 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_156_179 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_137_382 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_164_190 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_98_85 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_98_74 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_3_351 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_406 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_439 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_428 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_417 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_154_80 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_121_783 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_94_634 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_93_144 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_66_358 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_35_712 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_81_339 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5820_ hold870/Z _5827_/A2 _5821_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_35_778 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5751_ _5778_/A1 _5776_/A3 _5776_/A4 _5754_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_97_2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_175_411 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4702_ _4718_/A1 _4702_/A2 _4702_/B hold478/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_5682_ _5682_/A1 _5692_/A2 _5682_/A3 _5683_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand3_1
X_7421_ _7421_/D _7901_/RN _7872_/CLK _7995_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
X_4633_ _7993_/I _4652_/A1 _4636_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_8_61 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_175_499 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_162_105 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xhold602 hold602/I _7712_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
X_7352_ _7352_/D _7961_/RN _7505_/CLK _7352_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffsnq_1
X_4564_ _4564_/A1 _6537_/A2 _4568_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_7283_ hold4/I _7517_/Q _7279_/B _7283_/B _7284_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai31_1
Xmax_cap343 hold2/Z _6553_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__buf_12
Xhold613 hold613/I _7429_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
Xmax_cap354 _7901_/RN _7877_/RN VDD VSS gf180mcu_fd_sc_mcu7t5v0__buf_20
Xhold635 hold635/I _6079_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
Xhold624 hold624/I _4494_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
X_6303_ _4454_/Z _6315_/A2 _6303_/B _7783_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_6234_ _6545_/A1 hold6/Z _6234_/B hold67/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
Xhold657 _7722_/Q hold657/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
XFILLER_89_428 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4495_ hold247/Z _4504_/A2 hold248/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
Xhold646 _7560_/Q hold646/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
Xhold679 _7692_/Q hold679/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
Xhold668 hold668/I _7700_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
X_6165_ _7719_/Q _6174_/A2 _6166_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_112_761 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_69_141 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_940 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_951 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_962 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_5116_ _5309_/A1 _3723_/I _5344_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_2
X_6096_ _4460_/Z _6106_/A2 _6096_/B hold656/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
XTAP_973 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_984 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_995 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_5047_ _5006_/B _5254_/A2 _5254_/A3 _5689_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand3_4
XFILLER_45_509 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_72_317 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_25_233 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_53_531 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6998_ _7823_/Q _7202_/A2 _7202_/B1 _7783_/Q _7759_/Q _7202_/C2 _7000_/A3 VDD VSS
+ gf180mcu_fd_sc_mcu7t5v0__aoi222_1
X_5949_ _4476_/I _5953_/A2 _5949_/B hold354/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_80_372 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_13_428 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_43_25 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_179_783 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_40_247 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_166_477 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_166_455 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_127_809 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_7619_ _7619_/D _7853_/RN _7722_/CLK _7619_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_181_425 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_153_127 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_138_179 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_107_511 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_150_812 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_122_514 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_107_566 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_107_588 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_4_19 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_1_800 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_161_171 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_103_783 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_387 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_124_83 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_124_72 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_75_144 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_90_114 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_84_43 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_17_712 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_29_561 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_29_583 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_44_531 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_17_70 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_177_709 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_140_82 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_140_71 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_261 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_250 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_31_236 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XPHY_294 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_283 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_272 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_117_308 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_157_499 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_99_704 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_141_812 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_125_352 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_180_480 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_113_547 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_98_247 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_3_170 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4280_ _4280_/A1 _4280_/A2 _4274_/Z _4279_/Z _4281_/A4 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand4_1
XFILLER_98_258 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_67_601 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_79_472 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_39_303 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_12_2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7970_ _7970_/D _7323_/Z _7972_/CLK _7970_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_82_637 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6921_ _7660_/Q _7194_/B1 _6959_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_23_704 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_35_542 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6852_ _7133_/S _6852_/A2 _6852_/B _7928_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_5803_ _5803_/A1 _5803_/A2 _5803_/A3 _5803_/A4 _5804_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand4_1
XFILLER_62_394 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_50_534 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3995_ _7859_/Q _6452_/A1 _5988_/A1 _7641_/Q _3995_/C _3999_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi221_4
X_6783_ _6879_/A1 _6783_/A2 _6793_/C VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_22_247 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5734_ _5778_/A1 _5733_/Z _5737_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_5665_ _5665_/A1 _5753_/B _5671_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_30_291 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_163_425 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_135_105 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7404_ _7404_/D input75/Z _7410_/CLK _7404_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
X_4616_ _6539_/A1 _4618_/A2 _4616_/B _7409_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_163_469 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5596_ _5448_/B _5596_/A2 _5661_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_135_138 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_7335_ _7335_/D _7290_/Z _4398_/I1 _7335_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
Xhold410 hold410/I _4814_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
Xhold421 _4738_/Z _7454_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
XFILLER_150_108 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4547_ hold259/Z _4548_/A2 _4548_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_132_812 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xhold432 hold432/I _7640_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
Xhold443 hold443/I _7882_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
Xhold454 hold454/I _7592_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
Xhold465 hold465/I hold465/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
X_7266_ _7266_/A1 _7266_/A2 _7267_/C VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
Xhold476 _7988_/I hold476/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
Xhold487 _7583_/Q hold487/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
XFILLER_116_396 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4478_ hold716/Z _4487_/A1 _4482_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_6217_ hold64/Z _6225_/A2 _6217_/B _7743_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
Xhold498 hold498/I _6138_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
X_7197_ _7536_/Q _7197_/A2 _6938_/I _7392_/Q _7198_/A4 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_6148_ hold84/Z _6157_/A2 hold85/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_131_399 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_770 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_38_25 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_781 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_792 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_57_144 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_57_133 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_6079_ _4460_/Z _6089_/A2 _6079_/B hold636/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_26_531 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1925 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1914 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1903 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_159_709 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1958 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1947 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1936 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_14_737 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1969 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_110_30 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_41_567 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_139_411 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_110_74 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_167_753 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_182_734 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_166_263 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_154_414 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_139_499 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_126_105 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_182_789 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_123_812 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_1_641 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_103_580 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_103_591 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_37_807 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_95_97 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_151_70 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_91_423 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_151_92 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_91_456 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_17_542 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_32_534 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3780_ _4291_/B _3780_/A2 _7962_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_9_763 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_173_712 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_145_425 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5450_ _5643_/A2 _5608_/B _5752_/B1 _4996_/Z _5450_/C _5461_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi221_1
XFILLER_8_262 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4401_ _7425_/Q _4334_/Z _4402_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_5381_ _5022_/B _5381_/A2 _5382_/A3 _5381_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__or3_1
XFILLER_132_108 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_114_812 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4332_ _4292_/B _3738_/Z _4291_/B _4382_/A2 _7411_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai22_1
X_7120_ _7860_/Q _6938_/I _7188_/A2 _7381_/Q _7121_/A4 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_5_73 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_7051_ _7793_/Q _7190_/A2 _7190_/C1 _7703_/Q _7053_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_99_567 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_87_707 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4263_ _4263_/A1 _4263_/A2 _4263_/A3 _4263_/A4 _4282_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor4_1
XFILLER_140_174 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6002_ _4481_/I _6004_/A2 _6002_/B _7642_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_79_280 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4194_ _4194_/A1 _4194_/A2 _4194_/A3 _4194_/A4 _4202_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand4_1
XFILLER_94_250 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_39_144 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_39_155 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_7953_ _7953_/D _7959_/RN _4411_/I1 _7953_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_27_339 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_6904_ _6955_/A4 _6941_/A1 _7202_/C2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_4
XFILLER_23_512 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_23_523 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_35_361 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7884_ _7884_/D _7900_/RN _7892_/CLK _7884_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
X_6835_ _7643_/Q _6890_/A2 _6665_/Z _7747_/Q _6835_/C _6849_/B1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi221_1
XFILLER_11_707 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6766_ _6766_/A1 _6766_/A2 _6766_/A3 _6766_/A4 _6777_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand4_1
XFILLER_11_718 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_23_567 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_50_375 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_3978_ _7875_/Q _6486_/A1 hold150/I _7568_/Q _3994_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_5717_ _5717_/A1 _5717_/A2 _5717_/A3 _5718_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor3_1
Xclkbuf_2_1__f_mgmt_gpio_in[4] clkbuf_0_mgmt_gpio_in[4]/Z _4398_/I1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_108_105 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6697_ _6697_/A1 _6697_/A2 _6697_/A3 _6698_/C VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand3_1
X_5648_ _5648_/A1 _5648_/A2 _5624_/B _5648_/B2 _5648_/C _5743_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi221_1
XFILLER_40_37 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_156_37 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_151_417 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_5579_ _5669_/A1 _5027_/Z _5579_/B _5710_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_124_609 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_105_812 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7318_ _7901_/RN _4334_/Z _7318_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_151_428 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
Xhold251 _7615_/Q hold251/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
Xhold262 hold262/I _7829_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
Xhold240 hold240/I _6485_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
X_7249_ _7519_/Q _7249_/A2 _7251_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_132_664 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_131_141 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xhold273 _7773_/Q hold273/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
Xhold295 hold295/I _7594_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
XFILLER_78_707 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xhold284 hold284/I _7844_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
XFILLER_49_35 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_131_152 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_172_69 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_86_751 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2401 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_85_283 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_73_412 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1700 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_164_2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1733 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1722 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1711 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_121_51 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_54_681 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1766 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1755 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1744 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_121_73 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_14_534 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1799 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1777 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1788 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_81_77 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_14_589 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_41_375 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_81_99 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_155_712 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_6_700 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_6_744 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_142_406 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_114_108 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_6_788 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_182_597 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_114_119 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_107_182 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_146_92 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_146_70 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_122_130 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_111_804 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_46_8 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_96_559 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_110_369 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_76_261 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_76_250 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xinput8 mask_rev_in[13] input8/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XFILLER_39_90 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_49_486 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_91_242 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4950_ _5069_/A2 _4930_/Z _5458_/C _5015_/B _5357_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XFILLER_91_286 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3901_ _3901_/A1 _3901_/A2 _3901_/A3 _3901_/A4 _3917_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand4_1
X_4881_ hold819/Z _4882_/A2 hold820/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_3832_ hold609/Z _3886_/A2 _6520_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_4
XFILLER_60_673 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6620_ _7001_/C _4331_/Z _6621_/A2 _6620_/B _7918_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai31_1
X_6551_ hold233/Z _6553_/A2 _6551_/B hold276/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_3763_ _7973_/Q _7411_/Q _3763_/B _3764_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_5502_ _5502_/A1 _5652_/A3 _5767_/A2 _5641_/A2 _5509_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand4_1
X_3694_ hold66/I _3694_/ZN VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_158_594 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6482_ hold299/Z _6485_/A2 hold300/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_5433_ _5062_/Z _5176_/B _5624_/B _5482_/B2 _5433_/C _5434_/A4 VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai221_1
Xoutput301 _3961_/Z serial_data_1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__buf_4
XFILLER_145_299 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_133_428 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5364_ _5669_/A1 _5608_/B _5573_/A1 _5292_/B _5732_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_1
Xoutput334 _7948_/Q wb_dat_o[30] VDD VSS gf180mcu_fd_sc_mcu7t5v0__buf_4
Xoutput312 _7488_/Q wb_dat_o[10] VDD VSS gf180mcu_fd_sc_mcu7t5v0__buf_4
Xoutput323 _7482_/Q wb_dat_o[20] VDD VSS gf180mcu_fd_sc_mcu7t5v0__buf_4
XFILLER_160_258 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_160_247 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4315_ hold959/Z _4309_/S _4319_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_7103_ _7835_/Q _7203_/A2 _7204_/B1 _7771_/Q _7105_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_102_804 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_5295_ _5392_/A1 _5392_/A2 _5376_/B _5297_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor3_1
XFILLER_113_141 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7034_ hold66/I _7201_/A2 _7196_/A2 _7889_/Q _7035_/A4 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_4246_ _7814_/Q _6367_/A1 _7285_/A1 _7960_/Q _4248_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_142_17 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_95_570 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4177_ _7372_/Q _4522_/A1 _4574_/A1 _7394_/Q _7404_/Q _4599_/A1 _4179_/A3 VDD VSS
+ gf180mcu_fd_sc_mcu7t5v0__aoi222_1
XFILLER_67_283 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_27_103 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_7936_ _7936_/D _7938_/RN _7938_/CLK _7936_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XTAP_1029 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1007 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1018 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_7867_ _7867_/D _7901_/RN _7869_/CLK _7867_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
X_6818_ _7820_/Q _6880_/A2 _6893_/C1 _7634_/Q _6819_/A4 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_11_515 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_7798_ _7798_/D _7875_/RN _7863_/CLK _7798_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffsnq_1
XFILLER_51_25 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_167_36 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_137_712 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6749_ _7801_/Q _6883_/A2 _6883_/B1 _7785_/Q _6752_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_164_531 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_137_778 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_136_266 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_124_406 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_3_714 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_151_247 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_104_174 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_104_141 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_78_515 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_58_250 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_74_732 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_58_261 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_46_456 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_46_467 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2253 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2242 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2231 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2220 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_132_83 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_92_32 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_73_286 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_34_629 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2286 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2275 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2264 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1541 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1530 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_61_459 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_2297 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_159_303 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1585 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1574 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1563 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1552 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_25_70 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_30_802 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_70 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_81 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_42_673 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_92 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_1596 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_174_339 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_128_734 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_6_530 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_41_91 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_170_534 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_155_597 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_143_759 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_115_428 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_6_585 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_142_258 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_142_247 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_69_526 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_5080_ _5392_/A1 _5005_/Z _5779_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_2
XFILLER_123_494 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_123_483 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_96_323 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4100_ _4100_/A1 _4100_/A2 _4100_/A3 _4100_/A4 _4105_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand4_1
XFILLER_96_389 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4031_ _7786_/Q _6299_/A1 hold194/I _7351_/Q _4231_/B1 _4418_/I1 _4032_/A2 VDD VSS
+ gf180mcu_fd_sc_mcu7t5v0__aoi222_1
XFILLER_77_570 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_2_63 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_49_283 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_64_242 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5982_ hold366/Z _5987_/A2 _5983_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_4933_ _4917_/Z _4919_/Z _5201_/B _4941_/C VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi21_4
X_7721_ _7721_/D _7853_/RN _7805_/CLK _7721_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_177_111 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_177_144 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4864_ hold402/Z _4867_/A2 hold403/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_7652_ _7652_/D _7938_/RN _7653_/CLK _7652_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffsnq_1
XFILLER_119_712 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_3815_ hold72/Z hold609/Z _6503_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_4
X_7583_ _7583_/D _7923_/RN _7735_/CLK _7583_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
X_6603_ _7913_/Q _6586_/B _6609_/A2 _6604_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand3_1
X_4795_ _7228_/I0 _7484_/Q _4795_/S _7484_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_3746_ input58/Z _7411_/Q _3763_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_146_531 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6534_ hold233/Z _6536_/A2 _6534_/B hold279/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_118_266 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6465_ hold296/Z _6468_/A2 hold297/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_146_586 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5416_ _3722_/I _5709_/A1 _5452_/C _5543_/C _5417_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor4_4
X_3677_ _7932_/Q _7003_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_161_556 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_6396_ _6549_/A1 _6400_/A2 _6396_/B _7827_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
Xoutput175 _3699_/ZN mgmt_gpio_oeb[13] VDD VSS gf180mcu_fd_sc_mcu7t5v0__buf_4
X_5347_ _5768_/A2 _5680_/B1 _5347_/B _5347_/C _5353_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi211_1
Xoutput186 _3689_/ZN mgmt_gpio_oeb[23] VDD VSS gf180mcu_fd_sc_mcu7t5v0__buf_4
XFILLER_0_706 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
Xoutput197 _3679_/ZN mgmt_gpio_oeb[33] VDD VSS gf180mcu_fd_sc_mcu7t5v0__buf_4
XFILLER_101_100 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5278_ _5292_/B _5724_/B _5363_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_101_144 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7017_ _7776_/Q _7200_/A2 _7200_/B1 _7864_/Q _7023_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_4229_ _7527_/Q _4868_/A1 _4893_/A1 _7537_/Q _4236_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_47_209 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_101_166 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_46_69 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_55_286 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_7919_ _7919_/D _7961_/RN _7940_/CLK _7919_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_24_673 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_11_301 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_8_806 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_7_305 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_127_2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_152_534 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_124_203 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_109_288 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_109_277 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_124_247 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_105_461 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_133_792 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_87_54 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_78_389 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_59_570 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_47_732 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_19_445 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_46_264 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2061 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2050 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_61_212 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2094 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2083 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2072 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_61_278 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_159_144 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1393 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1382 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1360 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1371 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_70_790 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_42_492 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_175_637 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_128_531 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_128_520 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
Xinput22 mask_rev_in[26] input22/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyb_1
Xinput11 mask_rev_in[16] input11/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyb_1
X_4580_ hold757/Z _4583_/A2 _4581_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_30_676 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_162_309 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xinput44 mgmt_gpio_in[17] input44/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XFILLER_155_350 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xinput55 mgmt_gpio_in[27] input55/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyb_1
Xinput33 mask_rev_in[7] input33/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyb_1
Xinput66 mgmt_gpio_in[37] _8009_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyc_1
XFILLER_171_810 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_155_383 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xhold817 _7725_/Q hold817/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
Xhold828 hold828/I _6145_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
Xinput88 spimemio_flash_io1_oeb input88/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyb_1
Xinput77 ser_tx input77/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyb_1
Xhold806 _7830_/Q hold806/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
Xinput99 wb_adr_i[13] input99/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_143_567 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6250_ _6539_/A1 _6264_/A2 _6250_/B _7758_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
Xhold839 _7396_/Q hold839/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
X_5201_ _5200_/B _5230_/A1 _5663_/A1 _5201_/B _5371_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai31_1
XFILLER_170_353 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6181_ _4460_/Z _6191_/A2 _6181_/B _7726_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_42_2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5132_ _3722_/I _5087_/C _5006_/B _5254_/A2 _5643_/B1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor4_4
XFILLER_85_805 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_5063_ _5006_/C _5616_/A1 _5563_/B2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_4
XFILLER_65_551 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4014_ input30/Z _4249_/A2 _4232_/A2 input7/Z _6401_/A1 _7834_/Q _4016_/A2 VDD VSS
+ gf180mcu_fd_sc_mcu7t5v0__aoi222_1
XFILLER_38_743 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_92_392 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_37_286 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_5965_ hold698/Z _5970_/A2 _5966_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_4916_ _3728_/I _5369_/B _5230_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_4
X_7704_ _7704_/D _7938_/RN _7736_/CLK _7704_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
X_5896_ _6547_/A1 _5902_/A2 _5896_/B hold454/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_21_621 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7635_ _7635_/D _7877_/RN _7852_/CLK _7635_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_21_632 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4847_ _4454_/Z _4847_/A2 _4847_/B _7508_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_33_492 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_21_698 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_165_169 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4778_ _4454_/Z _4778_/A2 _4778_/B _7475_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_7566_ _7566_/D _7875_/RN _7567_/CLK _7566_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
X_3729_ _5369_/B _5022_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_8
XFILLER_134_523 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_106_203 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6517_ hold233/Z _6519_/A2 _6517_/B hold282/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_7497_ _7497_/D _7503_/CLK _7497_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_6448_ hold401/Z _6451_/A2 _6449_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_134_534 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_106_247 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_164_37 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6379_ _4476_/I _6383_/A2 _6379_/B hold238/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_115_770 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_88_676 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_90_318 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_71_510 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_28_275 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_29_798 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_44_702 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_113_96 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_43_223 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_157_659 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_156_103 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_12_676 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_153_810 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_137_350 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_138_93 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_180_673 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_113_707 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_78_120 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_429 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_418 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_407 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_94_602 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_120_250 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_66_315 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_93_156 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_74_392 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_19_286 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_5750_ _5754_/A1 _5754_/A2 _5775_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_175_401 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4701_ hold92/Z _3819_/Z _4701_/B _4702_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_5681_ _5681_/A1 _5620_/B _5681_/B _5723_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
XTAP_1190 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_4632_ _4652_/A1 _4632_/A2 _4632_/B hold574/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_7420_ _7420_/D _7901_/RN _7872_/CLK _7994_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_147_158 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_175_489 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
Xhold603 _7810_/Q hold603/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
X_7351_ _7351_/D _7961_/RN _7627_/CLK _7351_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffsnq_1
X_4563_ _4454_/Z _4563_/A2 _4563_/B _7388_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_7282_ _7282_/A1 _7282_/A2 _7282_/B _7283_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
Xmax_cap344 hold233/Z _4481_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__buf_12
XFILLER_116_534 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xhold636 hold636/I _7678_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
Xhold614 _7351_/Q hold614/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
Xhold625 hold625/I _7357_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
X_4494_ _4460_/Z _4504_/A2 _4494_/B hold625/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_6302_ hold871/Z _6315_/A2 _6303_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_6233_ hold66/Z hold6/Z _6234_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
Xhold669 _7864_/Q hold669/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
Xmax_cap355 _7875_/RN _7901_/RN VDD VSS gf180mcu_fd_sc_mcu7t5v0__buf_20
Xhold647 _7567_/Q hold647/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
Xhold658 _7626_/Q hold658/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
X_6164_ _4460_/Z _6174_/A2 _6164_/B _7718_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_112_751 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_85_602 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_930 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_941 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_952 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_58_805 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_5115_ _4999_/Z _5115_/A2 _5474_/B _5361_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_6095_ hold654/Z _6106_/A2 hold655/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_963 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_974 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_985 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_996 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_5046_ _5709_/A1 _5005_/Z _5404_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_111_283 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_150_28 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_65_392 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_25_212 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_53_521 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6997_ _6997_/A1 _6997_/A2 _6997_/A3 _6997_/A4 _6997_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__and4_1
X_5948_ hold353/Z _5953_/A2 _5949_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_178_250 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_178_283 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_166_412 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5879_ hold482/Z _5880_/A2 _5880_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_21_473 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_154_607 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7618_ _7618_/D _7923_/RN _7815_/CLK _7618_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_175_25 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_153_117 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_4_105 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7549_ _7549_/D _7308_/Z _4418_/I1 _7549_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffnrnq_1
XFILLER_153_139 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_147_692 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_4_116 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_162_673 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_134_364 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_68_34 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_68_45 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_1_812 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_103_762 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_76_602 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_333 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_102_250 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_88_495 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_48_304 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_75_134 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_90_104 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_75_156 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_91_638 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_56_392 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_16_256 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_31_215 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_251 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_240 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_169_283 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_157_434 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_295 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_284 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_273 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_262 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_129_103 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_33_70 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_157_489 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_126_810 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_98_204 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_152_183 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_4_672 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_79_451 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_140_389 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_121_570 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_94_421 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_82_605 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_66_167 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_54_307 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_54_318 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6920_ _6953_/A1 _6953_/A2 _6941_/A2 _7194_/B1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor3_4
X_6851_ _7928_/Q _7133_/S _6852_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_5802_ _5802_/A1 _5802_/A2 _5806_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_6782_ _7737_/Q _6878_/A2 _6783_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_3994_ _3994_/A1 _3994_/A2 _3994_/A3 _3995_/C VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand3_2
X_5733_ _5733_/A1 _5733_/A2 _5733_/A3 _5733_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__and3_1
XFILLER_175_242 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_148_467 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5664_ _5752_/B1 _5774_/A2 _5774_/B1 _5774_/A1 _5753_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_175_286 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5595_ _5661_/A1 _5662_/A1 _5319_/C _5596_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor3_1
Xclkbuf_leaf_54_csclk clkbuf_3_6__f_csclk/Z _7735_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
X_7403_ _7403_/D input75/Z _7410_/CLK _7403_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
X_4615_ hold763/Z _4618_/A2 _4616_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_4546_ hold233/Z _4548_/A2 _4546_/B _7381_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_7334_ _7334_/D _4440_/Z _4415_/A2 _7334_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
Xhold411 hold411/I _7494_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
Xhold400 hold400/I _7527_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
XFILLER_145_17 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_144_673 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_144_662 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
Xhold422 _7616_/Q hold422/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
XFILLER_116_342 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xhold433 _7802_/Q hold433/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
Xhold444 _7834_/Q hold444/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
Xhold466 hold466/I _7427_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
X_7265_ _7518_/Q _7265_/A2 _7265_/B1 _7519_/Q _7266_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_1
Xhold477 hold477/I _4702_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
XFILLER_131_312 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_89_215 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4477_ _4487_/A1 _6549_/A1 _4477_/B _7352_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
Xhold455 _7448_/Q hold455/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
X_6216_ hold68/Z _6225_/A2 _6217_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
Xhold488 _7716_/Q hold488/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
Xclkbuf_leaf_69_csclk _7528_/CLK _7649_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
X_7196_ _7547_/Q _7196_/A2 _7196_/B1 _7475_/Q _7198_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_1
Xhold499 hold499/I _7706_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
X_6147_ _4460_/Z _6157_/A2 _6147_/B hold577/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
XTAP_760 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_58_602 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_100_743 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_100_732 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_97_281 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_771 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_782 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_38_37 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_793 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_57_123 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_85_465 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6078_ hold634/Z _6089_/A2 hold635/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_5029_ _5643_/A2 _5027_/Z _5585_/B _5038_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_73_638 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_72_126 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_1915 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1904 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_81_660 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_38_392 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_54_25 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1959 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1948 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1937 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1926 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_81_671 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_13_215 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_14_727 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_54_69 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_179_570 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_110_64 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_182_702 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_21_281 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_181_212 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_154_459 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_5_425 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_119_73 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_162_481 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_122_345 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_79_99 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_150_676 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_122_389 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_103_570 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_49_602 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_174 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_64_605 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_36_318 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_49_668 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_151_60 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_91_446 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_76_487 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_48_189 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_151_82 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_32_502 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_71_170 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_9_753 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_172_212 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_157_286 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_117_128 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_4400_ _7430_/Q input77/Z _4400_/S _4400_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_5380_ _5380_/I _5641_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_126_673 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_126_662 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4331_ _7918_/Q _7575_/Q _7580_/Q _4331_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_140_142 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7050_ _7841_/Q _7204_/A2 _7204_/B1 _7769_/Q _7053_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_4262_ _4262_/A1 _4262_/A2 _4262_/A3 _4262_/A4 _4263_/A4 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand4_1
XFILLER_141_698 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_140_153 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_113_378 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6001_ hold660/Z _6004_/A2 _6002_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_4193_ input53/Z _5886_/A1 _4759_/A1 _7469_/Q _4194_/A4 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_7952_ _7952_/D _7959_/RN _4411_/I1 _7952_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_82_435 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_27_329 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_55_638 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_55_649 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6903_ _6908_/A1 _7913_/Q _6936_/A1 _6941_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand3_4
X_7883_ _7883_/D _7901_/RN _7899_/CLK _7883_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_35_373 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_6834_ _6834_/A1 _6834_/A2 _6834_/A3 _6834_/A4 _6835_/C VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand4_1
XFILLER_62_181 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_50_321 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6765_ hold57/I _6644_/Z _6665_/Z _7744_/Q _6891_/C1 _7778_/Q _6766_/A4 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi222_1
X_3977_ _7787_/Q _6299_/A1 _4219_/A2 input17/Z _3994_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_5716_ _5716_/A1 _5716_/A2 _5716_/A3 _5732_/A3 _5717_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand4_1
XFILLER_50_387 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6696_ _7847_/Q _6890_/B1 _6894_/C1 _7831_/Q _6697_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_163_234 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_163_212 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_136_459 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5647_ _4993_/B _5647_/A2 _5741_/A3 _5647_/B _5648_/C VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai31_1
X_5578_ _5578_/A1 _5578_/A2 _5578_/A3 _5578_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__and3_1
Xhold230 hold230/I _4685_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
X_7317_ _7901_/RN _4334_/Z _7317_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__and2_1
Xhold252 _7765_/Q hold252/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
Xhold241 hold241/I _7869_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
XFILLER_104_323 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4529_ _6539_/A1 _4531_/A2 _4529_/B _7373_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_7248_ _7248_/A1 _7277_/B _7248_/B _7951_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi21_1
Xhold263 _7465_/Q hold263/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
Xhold296 _7860_/Q hold296/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
Xhold285 _7366_/Q hold285/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
Xhold274 _7900_/Q hold274/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
XFILLER_172_37 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_132_676 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_131_164 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_104_389 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_105_31 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7179_ _7393_/Q _7200_/A2 _7201_/B1 _7507_/Q _7200_/B1 _7387_/Q _7182_/A1 VDD VSS
+ gf180mcu_fd_sc_mcu7t5v0__aoi222_1
XFILLER_86_763 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_85_240 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_590 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_46_605 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2402 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_18_318 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_45_104 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1734 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1723 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1712 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_121_41 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1701 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_157_2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1767 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1756 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1745 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1778 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1789 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_41_354 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_167_540 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_154_212 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_139_286 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_127_437 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_154_267 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_142_418 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_108_673 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_123_665 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_122_142 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_92_744 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xinput9 mask_rev_in[14] input9/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XFILLER_36_115 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_37_638 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_91_232 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_92_788 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_17_373 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3900_ _7813_/Q _6350_/A1 _6316_/A1 _7797_/Q _3901_/A4 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_60_630 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4880_ _6539_/A1 _4882_/A2 _4880_/B hold737/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_32_321 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3831_ hold26/Z hold41/Z hold75/Z _3963_/A4 _3886_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand4_4
X_3762_ _3762_/A1 _3762_/A2 _7974_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_6550_ hold274/Z _6553_/A2 hold275/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_20_538 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5501_ _5064_/B _5501_/A2 _5501_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__or2_1
XFILLER_72_2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_9_550 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_3693_ _7378_/Q _3693_/ZN VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_145_212 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6481_ _6549_/A1 _6485_/A2 _6481_/B _7867_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_5432_ _5778_/A1 _5162_/C _5686_/A2 _5725_/A1 _5435_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand4_1
XFILLER_161_738 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_105_109 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_5363_ _5600_/A1 _5363_/A2 _5797_/A1 _5363_/B _5703_/C VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai31_1
Xoutput335 _7949_/Q wb_dat_o[31] VDD VSS gf180mcu_fd_sc_mcu7t5v0__buf_4
Xoutput324 _7483_/Q wb_dat_o[21] VDD VSS gf180mcu_fd_sc_mcu7t5v0__buf_4
Xoutput302 _3927_/Z serial_data_2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__buf_4
Xoutput313 _7489_/Q wb_dat_o[11] VDD VSS gf180mcu_fd_sc_mcu7t5v0__buf_4
X_4314_ _4309_/S _4314_/A2 _4314_/B _7339_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_7102_ _7827_/Q _7202_/A2 _7202_/B1 _7787_/Q _7763_/Q _7202_/C2 _7105_/A2 VDD VSS
+ gf180mcu_fd_sc_mcu7t5v0__aoi222_1
XFILLER_99_354 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5294_ _5212_/Z _5294_/A2 _5294_/B _5299_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_114_676 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_141_495 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7033_ _7695_/Q _7194_/A2 _7202_/B1 _7785_/Q _7035_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_4245_ _7724_/Q hold28/I _4594_/A1 _7401_/Q _4858_/A1 _7523_/Q _4248_/A2 VDD VSS
+ gf180mcu_fd_sc_mcu7t5v0__aoi222_2
XFILLER_28_605 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4176_ _7605_/Q _5920_/A1 _4219_/A2 input12/Z _4176_/C _4179_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi221_1
XFILLER_67_273 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7935_ _7935_/D _7938_/RN _7935_/CLK _7935_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_24_811 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1008 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1019 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_7866_ _7866_/D _7901_/RN _7866_/CLK _7866_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_51_641 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_23_354 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6817_ _7682_/Q _6887_/B1 _6891_/B1 _7674_/Q _6819_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_7797_ _7797_/D _7853_/RN _7853_/CLK _7797_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_23_398 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6748_ _7639_/Q _6890_/A2 _6665_/Z hold68/I _6748_/C _6754_/B1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi221_1
XFILLER_50_195 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_176_392 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_129_6 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6679_ _7612_/Q _6647_/Z _6893_/B1 _7766_/Q _6681_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_136_256 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_152_738 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_151_215 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_117_481 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_2_247 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_120_602 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_104_164 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_78_527 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_116_63 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_76_34 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_19_638 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2210 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_100_392 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_74_744 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_73_221 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2243 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2232 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2221 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_46_479 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2287 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2276 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2265 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2254 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1542 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1531 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1520 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_92_77 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_61_438 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_14_321 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_27_682 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2298 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1575 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1564 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1553 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_60 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_71 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_82 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_175_808 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1597 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1586 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_41_151 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_93 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_174_318 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_167_381 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_127_212 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_143_716 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_10_593 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_41_70 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_182_384 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_170_524 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_157_70 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_170_579 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_110_156 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4030_ _4030_/A1 _4030_/A2 _4030_/A3 _4030_/A4 _4036_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand4_1
XFILLER_110_167 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_37_413 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_49_295 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5981_ hold16/Z _5987_/A2 _5981_/B hold17/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_64_276 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4932_ _4906_/S _5210_/B _5138_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_7720_ _7720_/D _7853_/RN _7720_/CLK _7720_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_80_747 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_52_449 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_178_602 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_17_192 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_32_140 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_33_641 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7651_ _7651_/D _7961_/RN _7960_/CLK _7651_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_178_646 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6602_ _6950_/A1 _6602_/A2 _7912_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_4863_ _4863_/A1 _7285_/A2 _4867_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_165_318 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3814_ hold53/Z hold37/Z _3843_/A3 _3864_/A4 hold609/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand4_4
XFILLER_119_702 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_4794_ _7227_/I0 _7483_/Q _4795_/S _7483_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_7582_ _7582_/D _7875_/RN _7830_/CLK _7582_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
X_3745_ _4292_/B _4284_/A1 _3745_/B _3747_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_158_392 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_119_724 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_118_212 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6533_ hold277/Z _6536_/A2 hold278/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_20_379 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_21_18 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_6464_ _6549_/A1 _6468_/A2 _6464_/B _7859_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_146_576 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5415_ _5415_/A1 _5415_/A2 _5415_/B _5521_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_133_215 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3676_ _7606_/Q _7027_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_133_248 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6395_ hold720/Z _6400_/A2 _6396_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
Xoutput176 _3698_/ZN mgmt_gpio_oeb[14] VDD VSS gf180mcu_fd_sc_mcu7t5v0__buf_4
X_5346_ _5692_/B _5692_/A2 _5347_/C VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_102_602 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xoutput198 _3678_/ZN mgmt_gpio_oeb[34] VDD VSS gf180mcu_fd_sc_mcu7t5v0__buf_4
Xoutput187 _3688_/ZN mgmt_gpio_oeb[24] VDD VSS gf180mcu_fd_sc_mcu7t5v0__buf_4
XFILLER_99_195 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_99_184 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_99_173 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5277_ _5624_/A1 _5431_/B _5566_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_7016_ _7016_/A1 _7016_/A2 _7016_/A3 _7016_/A4 _7026_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand4_1
XFILLER_87_357 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4228_ _7708_/Q _6141_/A1 _4759_/A1 _7468_/Q _4236_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_83_530 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_46_37 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4159_ _7621_/Q _5954_/A1 _4769_/A1 _7473_/Q _5971_/A1 _7629_/Q _4162_/A1 VDD VSS
+ gf180mcu_fd_sc_mcu7t5v0__aoi222_1
XFILLER_55_210 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_55_232 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_56_744 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_56_788 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_102_32 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_43_438 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_43_449 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7918_ _7918_/D _7961_/RN _7940_/CLK _7918_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_178_14 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_168_112 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7849_ _7849_/D _7877_/RN _7849_/CLK _7849_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_156_318 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_11_357 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_156_329 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_137_521 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_109_201 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_11_73 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_127_73 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_124_259 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_79_803 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_3_567 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_3_556 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_2_2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_78_368 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_47_722 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_19_424 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_46_210 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_46_254 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_46_276 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_47_799 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2051 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2040 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_62_747 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_159_101 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_2095 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2084 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2073 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2062 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1350 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_15_641 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_1383 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1361 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1372 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_30_600 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_42_460 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_159_156 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1394 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_14_195 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
Xinput12 mask_rev_in[17] input12/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyb_1
Xinput45 mgmt_gpio_in[18] input45/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyb_1
Xinput23 mask_rev_in[27] input23/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyb_1
Xinput34 mask_rev_in[8] input34/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyb_1
Xhold807 _7717_/Q hold807/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
Xinput56 mgmt_gpio_in[28] input56/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XFILLER_115_215 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xinput89 spimemio_flash_io2_do input89/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyb_1
Xinput78 spi_csb input78/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyb_1
Xhold818 _7510_/Q hold818/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
Xinput67 mgmt_gpio_in[3] input67/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_170_321 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_170_332 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xhold829 hold829/I _7709_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
XFILLER_115_248 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_115_237 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5200_ _5230_/A1 _5663_/A1 _5200_/B _5202_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_6180_ hold571/Z _6191_/A2 _6181_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_131_708 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_124_760 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5131_ _5006_/B _5344_/A2 _5480_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_69_335 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_35_2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_123_292 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5062_ _5006_/C _5616_/A1 _5062_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__and2_2
XFILLER_69_357 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4013_ _4013_/A1 _4013_/A2 _4013_/A3 _4013_/A4 _4013_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__and4_1
XFILLER_37_210 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_38_733 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_65_574 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_80_544 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_80_511 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_178_410 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7703_ _7703_/D _7923_/RN _7735_/CLK _7703_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
X_5964_ _6547_/A1 _5970_/A2 _5964_/B _7624_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_52_246 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_52_268 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4915_ _3728_/I _5369_/B _4915_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__and2_4
X_5895_ hold452/Z _5902_/A2 hold453/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_61_780 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_21_611 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_166_605 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7634_ _7634_/D _7877_/RN _7747_/CLK _7634_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_139_808 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4846_ hold824/Z _4847_/A2 _4847_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_138_318 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7565_ _7565_/D input75/Z _7567_/CLK _7565_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
X_6516_ hold280/Z _6519_/A2 hold281/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_20_176 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4777_ hold868/Z _4778_/A2 _4778_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_3728_ _3728_/I _5338_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_8
X_7496_ _7496_/D _7503_/CLK _7496_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_3659_ _5195_/B _5011_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_2
X_6447_ _6549_/A1 _6451_/A2 _6447_/B _7851_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_161_354 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6378_ hold237/Z _6383_/A2 _6379_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_5329_ _5431_/B _5624_/A2 _5540_/C _5335_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_114_270 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_559 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_180_37 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_29_700 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_29_722 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_180_59 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_91_809 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_56_530 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_16_405 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_44_747 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_31_408 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_169_443 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_24_460 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_157_649 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_156_115 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_137_340 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_8_659 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_152_321 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_152_365 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_98_76 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_419 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_408 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_94_636 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_78_176 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_19_265 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_47_91 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_47_574 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_170_70 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_62_522 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_19_298 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_179_229 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_34_246 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_43_780 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_148_605 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4700_ _3819_/Z hold64/I _4701_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_5680_ _5680_/A1 _5779_/A2 _5680_/B1 _5680_/B2 _5680_/C _5681_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi221_1
XTAP_1191 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1180 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_175_435 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4631_ hold34/Z _3830_/Z _4631_/B _4632_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_30_463 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_147_148 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7350_ _7350_/D _7961_/RN _7627_/CLK _7350_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffsnq_1
X_4562_ hold832/Z _4563_/A2 _4563_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_7281_ _7520_/Q _7281_/A2 _7281_/B1 _7518_/Q _7519_/Q _7281_/C2 _7282_/A2 VDD VSS
+ gf180mcu_fd_sc_mcu7t5v0__aoi222_1
XFILLER_171_641 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xhold615 _7597_/Q hold615/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
Xhold626 _7816_/Q hold626/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
X_4493_ hold623/Z _4504_/A2 hold624/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
Xhold604 _7529_/Q hold604/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
X_6301_ _6539_/A1 _6315_/A2 _6301_/B _7782_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_6232_ _4460_/Z hold6/Z _6232_/B _7750_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
Xmax_cap345 _4476_/I _6549_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__buf_8
XFILLER_143_354 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_89_419 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xhold659 _7650_/Q hold659/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
Xhold648 _7349_/Q hold648/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
Xhold637 _7579_/Q hold637/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
Xmax_cap356 _7875_/RN _7900_/RN VDD VSS gf180mcu_fd_sc_mcu7t5v0__buf_16
XFILLER_134_19 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6163_ hold630/Z _6174_/A2 _6164_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_920 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_931 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_942 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_953 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_5114_ _5648_/A1 _5058_/Z _5114_/A3 _5778_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand3_2
X_6094_ _4454_/Z _6106_/A2 _6094_/B hold921/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
XTAP_964 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_975 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_986 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_57_327 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5045_ _5538_/A1 _5042_/Z _5476_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_2
XFILLER_97_496 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_997 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_84_179 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_27_28 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_26_747 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_25_235 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6996_ _7669_/Q _7201_/B1 _7205_/A2 _7733_/Q _6997_/A4 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_5947_ _6547_/A1 _5953_/A2 _5947_/B _7616_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_139_627 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_5878_ _4454_/Z _5880_/A2 _5878_/B _7584_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_7617_ _7617_/D _7853_/RN _7805_/CLK _7617_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
X_4829_ _7503_/Q _4828_/S _4830_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_147_682 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_135_800 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_119_373 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7548_ _7548_/D _7307_/Z _4418_/I1 _7548_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffnrnq_1
XFILLER_146_170 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_134_321 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_107_546 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7479_ _7479_/D _7949_/CLK _7479_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_107_557 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_134_398 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_108_97 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_88_463 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_356 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_76_636 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_124_85 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_84_34 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_29_585 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_44_566 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_16_268 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_252 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_241 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_230 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_71_396 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_25_791 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_285 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_274 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_263 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_12_463 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_8_401 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_169_295 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_296 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_129_126 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_172_416 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_157_479 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_149_82 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_153_641 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_125_310 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_180_460 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_152_140 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_125_354 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_165_70 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_152_173 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_94_411 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_79_485 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_67_603 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xhold1 hold1/I hold1/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
XFILLER_66_179 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6850_ _7433_/Q _7927_/Q _6850_/B _6852_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_5801_ _5801_/A1 _5801_/A2 _5802_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_6781_ _7133_/S _6781_/A2 _6781_/B _7925_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_3993_ _7689_/Q _6090_/A1 _5971_/A1 _7633_/Q _3993_/C _3999_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi221_4
X_5732_ _5732_/A1 _5732_/A2 _5732_/A3 _5732_/A4 _5795_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand4_1
XFILLER_176_744 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5663_ _5663_/A1 _5753_/A2 _5774_/B1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_31_783 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_31_794 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_176_788 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_135_107 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5594_ _4969_/C _5606_/B _5599_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_4614_ _4614_/A1 _6537_/A2 _4618_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_7402_ _7402_/D input75/Z _7637_/CLK _7402_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
X_4545_ hold386/Z _4548_/A2 _4546_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
Xhold401 _7852_/Q hold401/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
XFILLER_135_129 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_129_682 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_7333_ _7901_/RN _4334_/Z _7333_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_116_321 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
Xhold434 _7866_/Q hold434/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
Xhold445 _7898_/Q hold445/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
Xhold423 _7786_/Q hold423/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
Xhold412 _7521_/Q hold412/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
X_7264_ _7520_/Q _7264_/A2 _7266_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
Xhold467 _7453_/Q hold467/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
Xhold478 hold478/I _7439_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
XFILLER_143_151 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4476_ _4476_/I _4750_/I1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_116_398 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xhold456 hold456/I _4729_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
Xhold489 _7806_/Q hold489/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
X_6215_ _4460_/Z _6225_/A2 _6215_/B _7742_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_131_357 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7195_ _7477_/Q _7195_/A2 _7195_/B1 _7471_/Q _7195_/C1 _7384_/Q _7198_/A2 VDD VSS
+ gf180mcu_fd_sc_mcu7t5v0__aoi222_1
X_6146_ hold575/Z _6157_/A2 hold576/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_750 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_761 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_100_722 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_772 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_783 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_794 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_100_788 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_85_477 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6077_ _4454_/Z _6089_/A2 _6077_/B hold760/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_57_168 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5028_ _5538_/A1 _5026_/Z _5545_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_85_499 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_85_488 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_72_105 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_38_371 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_38_360 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1916 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1905 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_53_330 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_54_37 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_159_6 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1949 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1938 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1927 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_14_717 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_41_525 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_53_352 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6979_ _7002_/B _6979_/A2 _6979_/A3 _6979_/B _7931_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai31_1
XFILLER_166_210 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_139_424 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_110_54 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_119_30 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_181_246 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_135_641 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_134_140 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_107_354 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_107_343 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_102_2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_79_34 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_162_460 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_79_89 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_135_73 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_89_783 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_142 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_49_658 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_95_99 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_91_425 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_29_371 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_48_179 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_56_190 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_60_812 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_158_766 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_158_744 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_157_243 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_157_221 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_13_783 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_157_298 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_173_769 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_172_257 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_181_780 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4330_ _4330_/I _7334_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_113_302 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_113_357 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_87_709 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4261_ _7347_/Q hold194/I _5988_/A1 _7636_/Q _4262_/A4 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_140_176 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_140_165 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6000_ _6549_/A1 _6004_/A2 _6000_/B _7641_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_140_187 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4192_ _7791_/Q _6316_/A1 _7285_/A1 _7961_/Q input21/Z _4239_/A2 _4194_/A3 VDD VSS
+ gf180mcu_fd_sc_mcu7t5v0__aoi222_1
XFILLER_95_753 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_28_809 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_7951_ _7951_/D _7959_/RN _4411_/I1 _7951_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_67_499 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_54_105 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7882_ _7882_/D _7900_/RN _7898_/CLK _7882_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_82_458 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6902_ _7912_/Q _7911_/Q _6936_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_4
XFILLER_54_138 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6833_ _7853_/Q _6890_/B1 _6894_/C1 _7837_/Q _6834_/A4 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_63_683 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_51_812 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_63_694 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_50_333 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_149_722 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_149_700 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_3976_ input40/Z _5903_/A1 hold43/I _7745_/Q _3996_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_6764_ _7379_/Q _6882_/A2 _6894_/C1 _7834_/Q _6764_/C _6766_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi221_1
XFILLER_11_709 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_148_210 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5715_ _5408_/C _5715_/A2 _5715_/A3 _5732_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor3_1
X_6695_ _7733_/Q _6830_/B _6889_/A2 _7701_/Q _6767_/C _6697_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi221_1
XFILLER_149_799 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_148_276 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_148_254 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5646_ _5510_/B _5646_/A2 _5646_/A3 _5740_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor3_1
XFILLER_164_747 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_163_224 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_40_39 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xhold220 hold220/I _5915_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
X_5577_ _5774_/A1 _4996_/Z _5062_/Z _5577_/B2 _5577_/C _5578_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi221_1
XFILLER_117_641 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_116_140 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_7316_ _7853_/RN _4334_/Z _7316_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__and2_1
Xhold231 hold231/I _7431_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
Xhold253 hold253/I _6264_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
Xhold242 _7861_/Q hold242/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
X_4528_ hold774/Z _4531_/A2 _4529_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_7247_ _7247_/A1 _7280_/A2 _7277_/B _7247_/C _7248_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi211_1
X_4459_ hold30/Z _3810_/S hold31/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
Xhold264 _4753_/Z _7465_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
Xhold275 hold275/I _6551_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
Xhold286 hold286/I _4513_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
Xhold297 hold297/I _6466_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
XFILLER_131_176 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_86_731 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7178_ _7178_/A1 _7178_/A2 _7178_/A3 _7184_/B1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor3_1
X_6129_ hold641/Z _6140_/A2 hold642/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_580 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_591 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_73_425 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_73_458 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_73_447 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1724 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1713 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_121_31 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1702 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_60_108 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_60_119 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_14_514 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_42_812 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1757 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1746 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1735 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_121_64 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_81_35 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_14_547 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_26_396 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1779 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1768 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_41_377 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_10_786 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_5_212 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_182_555 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_108_630 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_170_739 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_163_780 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_123_633 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_69_709 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_150_463 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_122_176 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_76_241 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_39_70 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_162_93 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_36_105 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_49_499 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xclkbuf_leaf_53_csclk clkbuf_3_6__f_csclk/Z _7597_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_33_812 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3830_ hold609/Z _3828_/I _3830_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__or2_4
Xclkbuf_leaf_68_csclk _7528_/CLK _7624_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
X_3761_ _7974_/Q _3752_/I _3762_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_5500_ _5064_/B _5501_/A2 _5641_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_158_585 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_146_747 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_145_224 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_118_449 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3692_ _7761_/Q _3692_/ZN VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_6480_ hold717/Z _6485_/A2 _6481_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_173_555 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5431_ _5624_/A1 _5648_/B2 _5431_/B _5625_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_65_2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_161_728 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5362_ _5362_/A1 _5520_/C _5362_/B1 _5362_/B2 _7539_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_126_460 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xoutput325 _7484_/Q wb_dat_o[22] VDD VSS gf180mcu_fd_sc_mcu7t5v0__buf_4
Xoutput303 _4414_/Z serial_load VDD VSS gf180mcu_fd_sc_mcu7t5v0__buf_4
Xoutput314 _7490_/Q wb_dat_o[12] VDD VSS gf180mcu_fd_sc_mcu7t5v0__buf_4
X_4313_ hold953/Z _4309_/S _4314_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_7101_ _7819_/Q _7207_/A2 _7207_/B1 _7721_/Q _7101_/C _7105_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi221_1
Xoutput336 _7499_/Q wb_dat_o[3] VDD VSS gf180mcu_fd_sc_mcu7t5v0__buf_4
X_7032_ _7687_/Q _7189_/B1 _7188_/A2 _7378_/Q _7035_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_5293_ _5561_/B _5293_/A2 _5293_/A3 _5293_/A4 _5298_/A4 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand4_1
XFILLER_113_176 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_101_327 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4244_ _7612_/Q _5937_/A1 _4853_/A1 _7521_/Q _4244_/C _4248_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi221_2
X_4175_ _7823_/Q _6384_/A1 _4614_/A1 _7410_/Q _4564_/A1 _7390_/Q _4179_/A1 VDD VSS
+ gf180mcu_fd_sc_mcu7t5v0__aoi222_1
XFILLER_83_712 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_55_425 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_83_778 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7934_ _7934_/D _7938_/RN _7935_/CLK _7934_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_42_108 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1009 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_7865_ _7865_/D _7900_/RN _7898_/CLK hold98/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_63_480 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_168_327 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7796_ _7796_/D _7923_/RN _7820_/CLK _7796_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
X_6816_ _7626_/Q _6659_/Z _6884_/B1 _7690_/Q _6819_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_23_344 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_168_349 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6747_ _6747_/A1 _6747_/A2 _6747_/A3 _6748_/C VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_149_563 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3959_ hold26/Z hold41/Z hold75/Z _3963_/A4 _3959_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__or4_2
XFILLER_164_511 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_6678_ _7732_/Q _6830_/B _6893_/C1 _7628_/Q _6767_/C _6681_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi221_1
X_5629_ _5079_/Z _5433_/C _5629_/B _5684_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_145_780 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_136_279 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_132_463 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_116_42 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_78_517 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_104_176 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_93_509 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_18_105 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_58_252 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2200 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_132_52 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_18_138 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2244 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2233 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2222 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2211 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_92_34 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_46_469 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2277 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2266 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2255 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1532 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1521 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1510 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_61_428 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2299 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2288 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_159_316 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1576 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1565 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1554 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1543 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_50 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_61 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_72 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_41_141 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_83 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_1598 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1587 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_14_388 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_94 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_128_747 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_182_352 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_182_330 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_6_543 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_127_279 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_108_460 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_151_761 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_123_441 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_173_70 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_151_783 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_150_282 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_123_496 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_96_347 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_110_179 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_65_712 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_92_531 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_37_425 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5980_ _7632_/Q _5987_/A2 _5981_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_65_778 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_24_108 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4931_ _5302_/A1 _5195_/B _5210_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__or2_1
XFILLER_52_439 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4862_ _4454_/Z _4862_/A2 _4862_/B hold888/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_7650_ _7650_/D _7961_/RN _7650_/CLK _7650_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
X_3813_ _3810_/S hold608/Z _3864_/A4 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_4
XFILLER_166_809 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6601_ _7912_/Q _6618_/A3 _6601_/B _6602_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_165_308 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4793_ _7226_/A1 _4795_/S _4793_/B _7482_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_20_325 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7581_ hold48/Z _7938_/RN _7606_/CLK _7581_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_32_185 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3744_ _3744_/A1 _3751_/A2 _4284_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_4
X_6532_ _6549_/A1 _6536_/A2 _6532_/B _7891_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_6463_ hold722/Z _6468_/A2 _6464_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_3675_ _7605_/Q _6707_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_134_717 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5414_ _5414_/A1 _5414_/A2 _5414_/A3 _5414_/A4 _5415_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor4_2
X_6394_ _6547_/A1 _6400_/A2 _6394_/B hold451/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
Xoutput177 _3697_/ZN mgmt_gpio_oeb[15] VDD VSS gf180mcu_fd_sc_mcu7t5v0__buf_4
X_5345_ _5176_/B _5573_/A1 _5477_/B2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_114_463 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_99_141 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_708 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xoutput199 _4393_/ZN mgmt_gpio_oeb[35] VDD VSS gf180mcu_fd_sc_mcu7t5v0__buf_4
Xoutput188 _3687_/ZN mgmt_gpio_oeb[25] VDD VSS gf180mcu_fd_sc_mcu7t5v0__buf_4
X_5276_ _5409_/B2 _5350_/A3 _5412_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_7015_ _7872_/Q _7195_/C1 _7015_/B _7016_/A4 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_4227_ _7668_/Q _6056_/A1 hold580/I _7571_/Q _4240_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_28_458 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4158_ _4158_/A1 _4158_/A2 _4158_/A3 _4158_/A4 _4204_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand4_2
XFILLER_56_734 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4089_ input54/Z _5886_/A1 _5971_/A1 _7630_/Q _4090_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_102_44 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_43_428 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7917_ _7917_/D _7961_/RN _7940_/CLK _7917_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_169_625 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_70_247 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_62_37 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_24_653 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_178_37 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7848_ _7848_/D _7877_/RN _7849_/CLK _7848_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffsnq_1
XFILLER_141_6 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_23_141 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_157_809 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_7779_ _7779_/D _7853_/RN _7877_/CLK _7779_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_168_179 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_164_341 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_109_235 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_180_812 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_164_396 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_152_558 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_87_34 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_87_12 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_160_591 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_133_783 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_105_496 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_78_325 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_47_712 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_143_84 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_143_73 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_101_691 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2052 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2041 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2030 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2085 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2074 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2063 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1340 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_61_236 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_15_653 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2096 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1384 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1362 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1373 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1351 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1395 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_174_105 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_128_522 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xinput13 mask_rev_in[18] input13/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyb_1
Xinput46 mgmt_gpio_in[19] input46/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyb_1
Xinput24 mask_rev_in[28] input24/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyb_1
Xinput35 mask_rev_in[9] input35/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XFILLER_171_812 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xinput57 mgmt_gpio_in[29] input57/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyb_1
Xhold808 _7584_/Q hold808/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
XFILLER_128_599 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_6_362 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
Xhold819 _7532_/Q hold819/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
Xinput79 spi_enabled _4396_/S VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
Xinput68 mgmt_gpio_in[5] input68/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyc_1
XFILLER_182_182 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_109_780 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5130_ _5735_/A2 _5179_/B _5749_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_5061_ _3722_/I _3723_/I _5006_/B _5616_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor3_4
XFILLER_28_2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_84_306 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4012_ _7712_/Q _6141_/A1 hold28/I _7728_/Q _4013_/A4 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_111_499 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_65_531 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
Xclkbuf_3_6__f_csclk clkbuf_0_csclk/Z clkbuf_3_6__f_csclk/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_80_534 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5963_ hold384/Z _5970_/A2 _5964_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_25_428 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4914_ _4914_/A1 _4914_/A2 _4914_/A3 _4914_/A4 _4914_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__or4_2
X_7702_ _7702_/D _7923_/RN _7737_/CLK _7702_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffsnq_1
X_5894_ _6545_/A1 _5902_/A2 hold96/Z hold97/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_7633_ _7633_/D _7877_/RN _7752_/CLK _7633_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
X_4845_ _6539_/A1 _4847_/A2 _4845_/B _7507_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_165_105 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7564_ _7564_/D input75/Z _7567_/CLK _7564_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffsnq_1
X_4776_ _6539_/A1 _4778_/A2 _4776_/B _7474_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_3727_ _3727_/I _5201_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__inv_8
X_6515_ _6549_/A1 _6519_/A2 _6515_/B _7883_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_20_199 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_180_108 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_162_812 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7495_ _7495_/D _7961_/RN _7876_/CLK _7495_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
X_3658_ _3658_/I _7282_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_134_525 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6446_ hold719/Z _6451_/A2 _6447_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_164_17 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6377_ _6547_/A1 _6383_/A2 _6377_/B _7818_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_5328_ _5333_/A3 _5495_/B2 _5540_/C VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_2
XFILLER_115_783 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_527 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_130_742 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_87_144 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_180_16 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5259_ _4996_/Z _5087_/B _5433_/C _5701_/C VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand3_2
XFILLER_29_712 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_83_394 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_28_277 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_71_567 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_169_499 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_156_127 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_156_105 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_132_2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_11_144 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_8_605 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_156_138 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_153_812 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_4_800 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_138_84 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_113_709 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_409 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_67_807 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_3_398 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_39_509 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_120_274 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_47_70 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_62_534 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_62_567 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1192 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1181 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1170 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_175_425 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4630_ _3830_/Z _4460_/Z _4631_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_175_447 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_8_53 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_162_108 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_144_812 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4561_ _6539_/A1 _4563_/A2 _4561_/B _7387_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_6300_ hold783/Z _6315_/A2 _6301_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_7280_ _4376_/B _7280_/A2 _7280_/A3 _7282_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand3_1
Xhold616 hold616/I _7437_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
Xhold627 _7694_/Q hold627/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
X_4492_ _4454_/Z _4504_/A2 _4492_/B hold900/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
Xhold605 hold605/I _4875_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
XFILLER_170_141 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6231_ hold563/Z hold6/Z _6232_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
Xmax_cap346 hold16/Z _6547_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_12
Xhold638 _7734_/Q hold638/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
Xhold649 _7367_/Q hold649/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
Xmax_cap357 _7938_/RN _7923_/RN VDD VSS gf180mcu_fd_sc_mcu7t5v0__buf_20
X_6162_ _4454_/Z _6174_/A2 _6162_/B _7717_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
XTAP_910 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_5113_ _5496_/A1 _5458_/C _5661_/A1 _5473_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor3_1
XFILLER_69_144 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_921 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_932 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_943 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_954 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_965 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_976 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_987 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_6093_ hold919/Z _6106_/A2 hold920/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_5044_ _5452_/C _5543_/C _5475_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_27_18 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_38_531 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_998 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_38_553 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_25_225 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_6995_ _7815_/Q _7207_/A2 _7207_/B1 _7717_/Q _7205_/B1 _7741_/Q _6997_/A3 VDD VSS
+ gf180mcu_fd_sc_mcu7t5v0__aoi222_1
XFILLER_53_567 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5946_ hold422/Z _5953_/A2 _5947_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_34_770 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_159_39 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5877_ hold808/Z _5880_/A2 _5878_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_166_414 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_138_105 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7616_ _7616_/D _7853_/RN _7811_/CLK _7616_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
X_4828_ _7228_/I0 _7502_/Q _4828_/S _7502_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_181_428 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_135_812 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4759_ _4759_/A1 _7285_/A2 _4763_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_7547_ _7547_/D _7875_/RN _7547_/CLK _7547_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_175_27 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7478_ _7478_/D _7949_/CLK _7478_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_161_141 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6429_ hold718/Z _6434_/A2 _6430_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_379 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_75_169 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_84_57 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_16_203 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_16_247 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_17_73 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_44_534 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_140_63 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_242 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_231 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_220 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_157_425 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_286 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_275 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_264 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_253 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_297 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_33_83 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_172_406 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_144_108 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_126_812 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_144_119 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_137_160 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_125_388 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_98_206 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_152_196 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_152_185 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_140_347 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_121_550 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_79_464 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
Xhold2 hold2/I hold2/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
XFILLER_181_70 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_94_478 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_63_810 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_47_372 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_47_383 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_5800_ _5800_/A1 _5800_/A2 _5801_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_3992_ _3992_/A1 _3992_/A2 _3992_/A3 _3993_/C VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand3_1
X_6780_ _7925_/Q _7133_/S _6781_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_90_673 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_35_567 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5731_ _5104_/B _5608_/B _5731_/B _5732_/A4 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_95_2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_175_222 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_148_447 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5662_ _5662_/A1 _5797_/A2 _5774_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_30_250 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_31_773 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_163_417 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_148_469 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5593_ _5608_/A1 _5167_/B _5606_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__or2_2
X_7401_ _7401_/D input75/Z _7401_/CLK _7401_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
X_4613_ _4454_/Z _4613_/A2 _4613_/B _7408_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_163_428 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7332_ _7901_/RN _4334_/Z _7332_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__and2_1
X_4544_ _6549_/A1 _4548_/A2 _4544_/B _7380_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_129_694 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
Xhold402 _7525_/Q hold402/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
X_7263_ _7263_/A1 _7277_/B _7263_/B _7954_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_144_664 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_143_141 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_132_804 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_128_193 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
Xhold435 hold435/I _6479_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
Xhold424 _8000_/I hold424/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
Xhold413 hold413/I _4855_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
X_4475_ hold216/Z hold49/Z _4475_/B hold217/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_4
Xhold468 hold468/I hold468/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
XFILLER_171_472 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6214_ hold695/Z _6225_/A2 _6215_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
Xhold446 hold446/I _6547_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
Xhold457 hold457/I _7448_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
Xhold479 _7572_/Q hold479/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
X_7194_ _7524_/Q _7194_/A2 _7194_/B1 _7505_/Q _7194_/C1 _7410_/Q _7199_/A2 VDD VSS
+ gf180mcu_fd_sc_mcu7t5v0__aoi222_1
X_6145_ _4454_/Z _6157_/A2 _6145_/B hold829/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
XTAP_740 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_751 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_97_283 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_97_294 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_85_423 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6076_ hold758/Z _6089_/A2 hold759/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_762 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_773 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_784 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_795 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_5027_ _5538_/A1 _5026_/Z _5027_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_85_467 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_85_445 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_166_8 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1906 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_26_534 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1939 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1928 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1917 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_6978_ _7604_/Q _6949_/I _6979_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_167_712 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_110_66 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5929_ hold539/Z _5936_/A2 hold540/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_179_594 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_139_447 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_110_99 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_70_59 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_70_37 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_22_784 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_182_726 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_126_108 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_108_801 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_21_283 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_182_737 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_119_171 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_119_42 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_150_601 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_1_611 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_110_509 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_95_209 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_88_250 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_95_45 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_95_89 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_95_67 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_45_810 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_151_73 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_72_673 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_17_567 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_32_504 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_157_233 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_12_250 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_145_428 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_138_480 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_172_247 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_126_664 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_114_804 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_153_483 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_125_141 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_4_460 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_153_494 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_140_133 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4260_ _4260_/A1 _4260_/A2 _4260_/A3 _4260_/A4 _4263_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand4_1
X_4191_ _7396_/Q _4579_/A1 _4774_/A1 _7475_/Q _4194_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_140_199 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_67_412 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_95_765 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_10_2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_7950_ _7950_/D _7959_/RN _7959_/CLK hold45/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_95_798 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_7881_ _7881_/D _7900_/RN _7881_/CLK _7881_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
X_6901_ _7931_/Q _7133_/S _6979_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_6832_ _7845_/Q _6894_/A2 _6659_/Z _7627_/Q _6834_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_51_802 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_149_712 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3975_ _7771_/Q _6265_/A1 _6418_/A1 _7843_/Q _3996_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_6763_ _6763_/A1 _6763_/A2 _6763_/A3 _6764_/C VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_176_531 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5714_ _5714_/A1 _5099_/B _5714_/B1 _5722_/A1 _5715_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai22_1
XFILLER_31_570 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_50_389 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6694_ _7839_/Q _6894_/A2 _6659_/Z _7621_/Q _6697_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_5645_ _5645_/A1 _5687_/B _5645_/A3 _5099_/B _5741_/A3 _5646_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai32_1
XFILLER_108_108 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_163_247 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5576_ _4960_/Z _5663_/A1 _5372_/Z _5576_/B2 _5576_/C _5715_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai221_1
Xhold210 _7707_/Q hold210/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
Xhold232 _7971_/Q hold232/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
Xhold221 hold221/I _7601_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
X_7315_ _7901_/RN _4334_/Z _7315_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__and2_1
Xhold243 hold243/I _6468_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
XFILLER_2_408 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4527_ _4527_/A1 _6537_/A2 _4531_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_4458_ hold49/Z hold387/Z _4461_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_7246_ _7246_/A1 _7246_/A2 _7247_/C VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_132_656 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
Xhold254 hold254/I _7765_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
XFILLER_116_196 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_104_347 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
Xhold265 _7885_/Q hold265/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
Xhold287 hold287/I _7366_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
Xhold276 hold276/I _7900_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
XFILLER_172_28 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_131_144 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
Xhold298 hold298/I _7860_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
X_7177_ _7177_/A1 _7177_/A2 _7177_/A3 _7177_/A4 _7178_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand4_1
XFILLER_105_33 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4389_ _4387_/S _7897_/Q _4389_/B _4389_/ZN VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
XTAP_570 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_6128_ _4454_/Z _6140_/A2 _6128_/B hold913/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_105_55 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_100_531 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_85_242 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_581 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_592 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_105_77 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_85_286 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6059_ hold910/Z _6072_/A2 _6060_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_58_478 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1725 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1714 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1703 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_53_150 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_54_673 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1758 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1747 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1736 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_81_481 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1769 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_167_564 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_127_428 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_154_247 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_6_747 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_107_141 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_123_645 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_122_122 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_122_100 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_107_196 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_1_441 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_89_570 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_103_380 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_1_496 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_92_724 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_77_798 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_91_212 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_64_459 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_36_139 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_55_70 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_72_492 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3760_ _3760_/A1 _3756_/B _3765_/A2 _3760_/B2 _7975_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_158_531 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_60_676 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_13_570 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_32_389 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_118_439 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3691_ _7769_/Q _3691_/ZN VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_5430_ _5247_/B _5724_/B _5550_/B _5725_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_173_567 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5361_ _5361_/A1 _5361_/A2 _5362_/B2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_1
Xoutput326 _7485_/Q wb_dat_o[23] VDD VSS gf180mcu_fd_sc_mcu7t5v0__buf_4
Xoutput304 _4413_/Z serial_resetn VDD VSS gf180mcu_fd_sc_mcu7t5v0__buf_4
Xoutput315 _7491_/Q wb_dat_o[13] VDD VSS gf180mcu_fd_sc_mcu7t5v0__buf_4
XFILLER_58_2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4312_ hold87/I _7414_/Q _4312_/B _4314_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_7100_ _7100_/A1 _7100_/A2 _7100_/A3 _7101_/C VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand3_1
X_5292_ _5724_/B _5624_/B _5292_/B _5293_/A4 VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
Xoutput337 _7500_/Q wb_dat_o[4] VDD VSS gf180mcu_fd_sc_mcu7t5v0__buf_4
XFILLER_113_144 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7031_ _7801_/Q _7191_/B1 _7194_/C1 _7809_/Q _7035_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_4243_ _4243_/A1 _4243_/A2 _4243_/A3 _4244_/C VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_19_19 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_68_743 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4174_ _4174_/A1 _4174_/A2 _4174_/A3 _4174_/A4 _4187_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand4_1
X_7933_ _7933_/D _7938_/RN _7938_/CLK _7933_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_67_286 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_36_673 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7864_ _7864_/D _7901_/RN _7864_/CLK _7864_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffsnq_1
X_7795_ _7795_/D _7853_/RN _7853_/CLK _7795_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
X_6815_ _6815_/A1 _6815_/A2 _6815_/A3 _6815_/A4 _6825_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand4_1
X_6746_ _7849_/Q _6890_/B1 _6894_/C1 _7833_/Q _6747_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_3958_ _3958_/A1 _4427_/B _3958_/B1 _3958_/B2 _7554_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_109_428 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3889_ _7627_/Q _5954_/A1 _4505_/A1 _7370_/Q _3892_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_6677_ _6677_/A1 _6677_/A2 _6677_/A3 _6677_/A4 _6684_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand4_1
XFILLER_164_534 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_164_556 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_136_247 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5628_ _5363_/B _5627_/Z _5634_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_5559_ _5559_/A1 _5415_/B _5560_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_2_205 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_104_166 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7229_ _7949_/Q _7228_/S _7230_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_104_199 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_76_58 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_86_562 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_59_798 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2201 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_73_234 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_73_212 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_18_128 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2234 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2223 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2212 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_132_75 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_92_24 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_2278 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2267 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2256 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2245 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_162_2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1533 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1522 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1511 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1500 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_40 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_42_621 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2289 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1566 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1555 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1544 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_51 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_62 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_73 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_1599 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1588 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1577 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_25_73 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_84 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_42_676 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_95 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_155_567 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_170_504 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_143_718 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_69_507 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_150_250 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_110_103 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_37_415 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_49_297 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_49_286 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_92_565 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_52_407 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_4930_ _5195_/B _5201_/B _5210_/A3 _4926_/Z _4930_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__or4_4
XFILLER_80_727 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_17_150 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4861_ hold886/Z _4862_/A2 hold887/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_3812_ hold607/Z _7342_/Q _7414_/Q _3812_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_6600_ _7434_/Q _6599_/Z _6601_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_4792_ _7482_/Q _4795_/S _4793_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_7580_ _7580_/D _7961_/RN _7624_/CLK _7580_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_2
X_3743_ _7346_/Q _7345_/Q _7344_/Q _4206_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor3_4
X_6531_ hold728/Z _6536_/A2 _6532_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_3674_ _7957_/Q _7278_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_146_534 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_118_247 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6462_ _6547_/A1 _6468_/A2 _6462_/B hold429/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_5413_ _5732_/A1 _5413_/A2 _5413_/A3 _5588_/A3 _5414_/A4 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand4_1
X_6393_ hold449/Z _6400_/A2 hold450/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_5344_ _5344_/A1 _5344_/A2 _5623_/A1 _5350_/A3 _5545_/A2 _5687_/B _5347_/B VDD VSS
+ gf180mcu_fd_sc_mcu7t5v0__oai33_1
Xoutput167 _4431_/Z debug_in VDD VSS gf180mcu_fd_sc_mcu7t5v0__buf_4
Xoutput178 _3696_/ZN mgmt_gpio_oeb[16] VDD VSS gf180mcu_fd_sc_mcu7t5v0__buf_4
Xoutput189 _3686_/ZN mgmt_gpio_oeb[26] VDD VSS gf180mcu_fd_sc_mcu7t5v0__buf_4
XFILLER_101_114 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_5275_ _5714_/B1 _5623_/A1 _5712_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_141_283 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7014_ _7014_/A1 _7014_/A2 _7015_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_4226_ _7558_/Q _5817_/A1 _4522_/A1 _7371_/Q _4267_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_4157_ _7661_/Q _6039_/A1 _6333_/A1 _7799_/Q _4158_/A4 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_95_381 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_83_532 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_46_28 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_46_39 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_55_212 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_55_223 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4088_ _7349_/Q hold194/I _4249_/A2 input26/Z _4505_/A1 _7365_/Q _4090_/A2 VDD VSS
+ gf180mcu_fd_sc_mcu7t5v0__aoi222_2
XFILLER_102_34 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_102_23 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7916_ _7916_/D _7923_/RN _7935_/CLK _7916_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_71_738 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_70_204 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7847_ _7847_/D _7875_/RN _7847_/CLK _7847_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffsnq_1
XFILLER_169_648 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_169_637 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_23_153 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_24_676 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_24_665 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_7778_ _7778_/D _7877_/RN _7851_/CLK _7778_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
X_6729_ _6729_/A1 _6729_/A2 _6729_/A3 _6728_/Z _6731_/B1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand4_1
XFILLER_164_353 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_137_567 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xclkbuf_leaf_52_csclk clkbuf_3_6__f_csclk/Z _7698_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_11_31 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_127_42 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_3_514 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_11_97 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_133_773 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_132_250 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_120_401 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_87_68 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_132_283 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_120_456 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_87_79 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
Xclkbuf_leaf_67_csclk clkbuf_3_3__f_csclk/Z _7653_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_120_467 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_143_96 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_86_392 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2042 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2020 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2031 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_62_727 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_61_226 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_61_215 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_15_621 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2086 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2075 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2064 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2053 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1341 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1330 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2097 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1363 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1374 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1352 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_30_602 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_42_473 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_1396 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1385 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_156_810 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_30_668 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_128_534 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xinput14 mask_rev_in[19] input14/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyb_1
Xinput25 mask_rev_in[29] input25/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyb_1
Xinput36 mgmt_gpio_in[0] input36/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyc_1
XFILLER_155_375 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_116_729 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
Xinput69 mgmt_gpio_in[6] input69/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XFILLER_10_392 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
Xhold809 _7522_/Q hold809/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
Xinput47 mgmt_gpio_in[1] input47/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyb_1
Xinput58 mgmt_gpio_in[2] input58/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__buf_3
XFILLER_143_559 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_124_751 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_97_602 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_170_389 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_151_570 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5060_ _5319_/C _5692_/B _5301_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_123_283 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_84_318 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4011_ _7736_/Q _6192_/A1 _6090_/A1 _7688_/Q _4013_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_77_392 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_37_212 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5962_ hold64/Z _5970_/A2 _5962_/B hold77/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_25_418 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_53_738 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4913_ _4914_/A1 _4914_/A2 _4914_/A3 _4914_/A4 _5211_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor4_4
X_7701_ _7701_/D _7938_/RN _7733_/CLK _7701_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffsnq_1
X_5893_ hold95/Z _5902_/A2 hold96/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_61_760 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_7632_ hold17/Z _7877_/RN _7747_/CLK _7632_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
X_4844_ hold752/Z _4847_/A2 _4845_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_7563_ _7563_/D _7875_/RN _7563_/CLK _7563_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
X_4775_ hold782/Z _4778_/A2 _4776_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_3726_ _5199_/B _5200_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__inv_8
X_6514_ hold721/Z _6519_/A2 _6515_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_146_342 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_134_504 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_119_567 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_107_718 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7494_ _7494_/D _7961_/RN _7572_/CLK _7494_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
X_6445_ hold16/Z _6451_/A2 hold60/Z hold61/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_3657_ _7916_/Q _6905_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_2
X_6376_ hold528/Z _6383_/A2 _6377_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_114_250 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_88_624 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_88_602 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5327_ _5431_/B _5624_/A2 _5803_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_506 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_102_423 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_102_467 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5258_ _5290_/B _5409_/B2 _5258_/B _5585_/C VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_5189_ _5658_/B _5643_/A2 _5642_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_68_392 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4209_ _4075_/B _3959_/Z hold580/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_113_55 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_113_44 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_28_256 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_43_215 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_43_237 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_12_602 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_52_771 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_12_646 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_125_2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_165_651 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_125_548 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_98_34 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_4_812 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_180_676 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_106_751 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_98_45 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_152_389 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_133_570 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_98_89 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_105_283 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_94_605 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_19_212 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_19_223 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_47_532 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_47_93 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_63_70 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_179_70 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1182 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1171 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1160 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_270 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_179_92 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_175_415 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_147_117 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_1193 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_4560_ hold750/Z _4563_/A2 _4561_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_30_498 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
Xhold617 _7438_/Q hold617/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
X_4491_ hold898/Z _4504_/A2 hold899/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
Xhold606 hold606/I _7529_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
Xmax_cap347 hold63/Z _6545_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__buf_12
X_6230_ _4454_/Z hold6/Z _6230_/B _7749_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_131_507 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xhold628 hold628/I _6113_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
Xhold639 hold639/I _6198_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
Xmax_cap358 input75/Z _7938_/RN VDD VSS gf180mcu_fd_sc_mcu7t5v0__buf_20
XFILLER_171_698 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_6161_ hold807/Z _6174_/A2 _6162_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_40_2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_900 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_5112_ _4996_/Z _5793_/A2 _5673_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_911 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_922 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_933 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_944 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_112_765 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6092_ hold47/Z _6106_/A2 _6092_/B hold622/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_69_156 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_955 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_966 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_977 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_5043_ _5548_/A1 _5043_/A2 _5543_/C VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_4
XFILLER_111_286 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_85_649 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_85_638 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_38_521 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_988 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_999 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
Xclkbuf_0_wbbd_sck _7958_/Q clkbuf_0_wbbd_sck/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_93_693 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_81_811 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_25_215 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_80_321 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6994_ _7879_/Q _7203_/B1 _7204_/A2 _7839_/Q _6997_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_5945_ hold64/I _5953_/A2 _5945_/B _7615_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_34_760 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5876_ _4460_/Z _5880_/A2 _5876_/B _7583_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_33_281 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7615_ _7615_/D _7853_/RN _7720_/CLK _7615_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffsnq_1
X_4827_ _7227_/I0 _7501_/Q _4828_/S _7501_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_166_459 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_138_128 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4758_ _4454_/Z _4758_/A2 _4758_/B _7467_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_7546_ _7546_/D _7875_/RN _7830_/CLK _7546_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_146_183 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4689_ hold367/Z _3819_/Z _4689_/B _4690_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_134_323 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3709_ _7631_/Q _3709_/ZN VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_4_108 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_7477_ _7477_/D input75/Z _7477_/CLK _7477_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
X_6428_ _6547_/A1 _6434_/A2 _6428_/B _7842_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_162_676 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_161_175 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_134_389 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_115_570 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6359_ hold603/Z _6366_/A2 _6360_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_115_581 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_68_37 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_314 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_103_776 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_88_476 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_76_605 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_130_595 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_103_798 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_88_487 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_76_638 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_48_318 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_124_98 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_90_129 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_90_118 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_29_565 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_17_749 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_140_75 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_210 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_31_207 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_243 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_232 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_221 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_71_398 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_276 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_265 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_254 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_169_297 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_169_286 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_298 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_287 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_33_73 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_149_73 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_153_665 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_99_708 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_180_484 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_152_164 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_4_664 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_3_141 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_140_326 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_79_421 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_79_410 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_121_540 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
Xhold3 hold3/I hold3/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
XFILLER_67_638 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_90_630 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_62_321 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3991_ _7665_/Q _6039_/A1 _6192_/A1 _7737_/Q _3992_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_23_708 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5730_ _5763_/A3 _5730_/A2 _5738_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_176_702 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_175_212 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5661_ _5661_/A1 _5661_/A2 _5661_/B _5774_/C VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_88_2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7400_ _7400_/D input75/Z _7477_/CLK _7400_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
X_5592_ _5608_/A1 _5167_/B _5753_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_4612_ hold836/Z _4613_/A2 _4613_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_7331_ _7901_/RN _4334_/Z _7331_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__and2_1
X_4543_ hold731/Z _4548_/A2 _4544_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_7262_ _7262_/A1 _7280_/A2 _7277_/B _7262_/C _7263_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi211_1
Xhold436 hold436/I _7866_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
Xhold425 hold425/I _5892_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
Xhold414 hold414/I _7521_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
Xhold403 hold403/I _4865_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
Xhold469 hold469/I _7419_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
X_4474_ hold49/Z _7268_/A1 _4475_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_144_676 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_143_175 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_143_153 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xhold458 _7873_/Q hold458/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
XFILLER_116_389 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xhold447 hold447/I _7898_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
X_6213_ _4454_/Z _6225_/A2 _6213_/B _7741_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_7193_ _7396_/Q _7193_/A2 _7193_/B1 _7473_/Q _7193_/C1 _7532_/Q _7199_/A1 VDD VSS
+ gf180mcu_fd_sc_mcu7t5v0__aoi222_1
X_6144_ hold827/Z _6157_/A2 hold828/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_730 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_741 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_752 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_58_605 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xload_slew350 hold5/Z _6537_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__buf_20
X_6075_ hold47/Z _6089_/A2 _6075_/B hold365/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
XTAP_763 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_774 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_785 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_5026_ _5548_/A1 _5535_/A1 _5026_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__and2_1
XTAP_796 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1907 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_81_641 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_54_17 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_54_39 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1929 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1918 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_53_354 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6977_ _7210_/A2 _6977_/A2 _6977_/A3 _6977_/A4 _6979_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor4_1
XFILLER_179_540 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_110_34 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5928_ hold64/I _5936_/A2 _5928_/B hold154/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_53_398 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_22_741 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_34_590 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_166_212 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5859_ _7576_/Q _5868_/A2 _5860_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_21_240 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_166_267 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_181_215 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_166_278 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_135_621 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_119_21 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_5_428 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7529_ _7529_/D _7938_/RN _7741_/CLK _7529_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_181_248 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_119_98 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_150_646 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_134_186 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_122_337 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_89_774 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_177 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_49_638 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_130_392 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_28_62 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_91_438 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_44_321 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_32_538 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_44_50 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_44_387 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_44_398 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_157_212 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_9_712 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_12_273 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_145_418 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_172_259 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_125_120 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_126_676 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_5_77 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_5_99 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4190_ _7783_/Q _6299_/A1 _6418_/A1 _7839_/Q _7580_/Q _5870_/A1 _4194_/A1 VDD VSS
+ gf180mcu_fd_sc_mcu7t5v0__aoi222_1
XFILLER_94_210 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_67_424 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_121_381 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_82_427 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7880_ _7880_/D _7901_/RN _7899_/CLK _7880_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffsnq_1
XFILLER_85_90 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_63_641 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6900_ _7133_/S _6900_/A2 _6900_/B _7930_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_35_310 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6831_ _7707_/Q _6889_/A2 _6834_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_90_460 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_35_354 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3974_ _7657_/Q _6022_/A1 _6367_/A1 _7819_/Q _3989_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_6762_ _7664_/Q _6885_/A2 _6893_/B1 _7770_/Q _6763_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_176_510 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_176_521 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_148_212 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5713_ _5716_/A1 _5716_/A2 _5716_/A3 _5795_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand3_1
X_6693_ _7613_/Q _6647_/Z _6887_/B1 _7677_/Q _6705_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_148_256 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5644_ _5644_/A1 _5644_/A2 _5644_/A3 _5804_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_163_215 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_156_19 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5575_ _5212_/Z _5575_/A2 _5768_/A3 _5576_/C VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand3_1
Xhold200 hold200/I _6123_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
Xhold211 hold211/I _6140_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
X_7314_ _7900_/RN _4334_/Z _7314_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_172_771 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xhold233 hold233/I hold233/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
Xhold222 _7713_/Q hold222/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
XFILLER_116_164 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xhold244 hold244/I _7861_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
X_4526_ _4454_/Z _4526_/A2 _4526_/B _7372_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_7245_ _7520_/Q _7245_/A2 _7245_/B1 _7519_/Q _7246_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_131_123 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_116_186 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
Xhold266 hold266/I _6519_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
Xhold255 _7893_/Q hold255/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
Xhold277 _7892_/Q hold277/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
X_4457_ hold648/Z _4487_/A1 _4462_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_49_17 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_132_668 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xhold288 _7828_/Q hold288/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
Xhold299 _7868_/Q hold299/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
X_7176_ _7391_/Q _6938_/I _7188_/A2 _7756_/Q _7177_/A4 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_105_23 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_4388_ _4387_/S input92/Z _4389_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_86_733 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_560 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_6127_ hold911/Z _6140_/A2 hold912/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_112_392 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_86_744 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_85_232 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_571 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_582 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_593 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_6058_ hold47/Z _6072_/A2 _6058_/B _7668_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_5009_ _5199_/B _4898_/Z _4915_/Z _5005_/Z _5529_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand4_4
XFILLER_26_321 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_39_682 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1715 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1704 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_53_140 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1748 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1737 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1726 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1759 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_41_357 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_139_212 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_10_744 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_182_524 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_155_738 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_108_632 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_108_676 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_146_52 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_135_484 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_122_112 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_146_85 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_150_487 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_110_318 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_39_50 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_49_424 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_39_61 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_76_254 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_18_800 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_92_747 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_91_246 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_17_354 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_45_641 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_60_611 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_55_82 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_177_318 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_32_346 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_44_184 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_13_560 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_71_70 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_145_215 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3690_ _7777_/Q _3690_/ZN VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_5360_ _5415_/B _5360_/A2 _5360_/B _7279_/B _5361_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_114_602 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xoutput305 _4430_/Z spi_sdi VDD VSS gf180mcu_fd_sc_mcu7t5v0__buf_4
Xoutput316 _7492_/Q wb_dat_o[14] VDD VSS gf180mcu_fd_sc_mcu7t5v0__buf_4
X_4311_ _7414_/Q _4308_/S _4311_/A3 _4312_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor3_1
X_5291_ _5624_/B _5759_/A1 _5431_/B _5292_/B _5291_/C _5293_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi221_1
Xoutput327 _7942_/Q wb_dat_o[24] VDD VSS gf180mcu_fd_sc_mcu7t5v0__buf_4
Xoutput338 _7501_/Q wb_dat_o[5] VDD VSS gf180mcu_fd_sc_mcu7t5v0__buf_4
XFILLER_113_156 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_99_357 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7030_ _7133_/S _7030_/A2 _7030_/B _7933_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_4242_ _7732_/Q _6192_/A1 _4589_/A1 _7399_/Q _4243_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_141_487 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_101_329 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4173_ _7709_/Q _6141_/A1 hold28/I _7725_/Q _4174_/A4 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_95_574 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7932_ _7932_/D _7938_/RN _7938_/CLK _7932_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_169_808 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_7863_ _7863_/D _7875_/RN _7863_/CLK _7863_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffsnq_1
XFILLER_168_318 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7794_ _7794_/D _7853_/RN _7853_/CLK _7794_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
X_6814_ _7754_/Q _6644_/Z _6665_/Z _7746_/Q _6891_/C1 _7780_/Q _6815_/A4 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi222_1
XFILLER_23_357 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_168_329 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6745_ _7735_/Q _6830_/B _6889_/A2 _7703_/Q _6767_/C _6747_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi221_1
XFILLER_11_519 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3957_ hold946/Z _4284_/A1 _4427_/B _3958_/B2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_137_705 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_50_176 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3888_ _7781_/Q _6282_/A1 _6418_/A1 _7845_/Q _3892_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_6676_ _7700_/Q _6889_/A2 _6890_/A2 _7636_/Q _6677_/A4 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_5627_ _5741_/B _5627_/A2 _5627_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__and2_1
X_5558_ _5542_/Z _5557_/Z _5558_/B _5640_/B1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_4509_ _4454_/Z _4521_/A2 _4509_/B hold909/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_5489_ _5548_/A1 _5150_/Z _5497_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_120_605 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7228_ _7228_/I0 _7948_/Q _7228_/S _7948_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_104_189 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_116_99 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_7159_ _7159_/A1 _7159_/A2 _7159_/A3 _7159_/A4 _7160_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__or4_1
XFILLER_76_37 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_59_766 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_390 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_74_747 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2235 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2224 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2213 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2202 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_132_65 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_27_641 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2268 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2257 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2246 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1523 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1512 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1501 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_92_69 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_30 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_54_482 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2279 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_159_307 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_155_2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1567 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1556 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1545 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1534 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_81_290 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_41 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_52 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_26_195 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_63 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_74 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_1589 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1578 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_85 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_96 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_128_727 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_127_215 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_182_332 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_157_51 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_127_237 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_6_534 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_6_523 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_41_73 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_157_73 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_155_579 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_143_708 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_136_771 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_182_387 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_170_538 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_111_638 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_2_784 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_110_148 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_1_283 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_2_34 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_37_438 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_80_717 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_65_769 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_64_246 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_73_780 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_33_600 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_178_605 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4860_ hold47/Z _4862_/A2 _4860_/B hold599/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_3811_ _3810_/S _3808_/Z _3811_/B _3843_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi21_4
XFILLER_60_463 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_6530_ _6547_/A1 _6536_/A2 _6530_/B hold440/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_32_176 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4791_ _7224_/I0 _7481_/Q _4795_/S _7481_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_3742_ _7346_/Q _7345_/Q _3751_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_2
XFILLER_70_2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3673_ _3673_/I _7273_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_6461_ hold427/Z _6468_/A2 hold428/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_173_354 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6392_ _6545_/A1 _6400_/A2 _6392_/B hold463/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_5412_ _5585_/A1 _5793_/A2 _5412_/B _5588_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_5343_ _5343_/A1 _5343_/A2 _5354_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_114_454 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_99_132 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xoutput168 _7982_/Z irq[0] VDD VSS gf180mcu_fd_sc_mcu7t5v0__buf_4
Xoutput179 _3695_/ZN mgmt_gpio_oeb[17] VDD VSS gf180mcu_fd_sc_mcu7t5v0__buf_4
XFILLER_102_605 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_101_104 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_87_305 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5274_ _5292_/B _5431_/B _5706_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_114_498 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7013_ _7896_/Q _7197_/A2 _6938_/I _7856_/Q _7014_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_4225_ _7790_/Q _6316_/A1 _4604_/A1 _7405_/Q _4267_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_4156_ _7767_/Q _6265_/A1 hold150/I _7564_/Q _4604_/A1 _7406_/Q _4158_/A3 VDD VSS
+ gf180mcu_fd_sc_mcu7t5v0__aoi222_2
XFILLER_68_585 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_28_449 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_56_747 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4087_ _7848_/Q _6435_/A1 _6384_/A1 _7824_/Q _4090_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_7915_ _7915_/D _7923_/RN _7938_/CLK _7915_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffsnq_2
XFILLER_36_460 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_63_290 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_62_17 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7846_ _7846_/D _7875_/RN _7847_/CLK _7846_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffsnq_1
X_4989_ _5006_/B _5006_/C _5344_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_4
X_7777_ _7777_/D _7901_/RN _7829_/CLK _7777_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_23_198 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_51_496 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_177_682 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_165_800 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_137_513 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_6728_ _6728_/A1 _6728_/A2 _6728_/A3 _6728_/A4 _6728_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__and4_1
XFILLER_164_321 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_109_215 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_6659_ _6878_/A2 _6665_/A2 _6659_/A3 _6659_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__and3_2
XFILLER_152_516 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_164_398 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_118_771 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_117_292 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_105_443 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_132_262 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_78_327 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_94_809 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_143_53 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_100_170 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_74_511 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2010 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_74_566 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2043 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2021 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2032 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_62_739 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_62_717 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_15_611 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_46_268 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_55_780 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2076 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2065 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2054 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1331 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1320 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2098 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2087 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1364 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1375 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1353 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1342 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_463 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1397 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1386 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_14_176 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_42_496 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_30_658 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_168_61 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
Xinput37 mgmt_gpio_in[10] input37/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyb_1
Xinput15 mask_rev_in[1] input15/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyb_1
Xinput26 mask_rev_in[2] input26/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XFILLER_155_354 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_155_343 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
Xinput59 mgmt_gpio_in[30] input59/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyc_1
Xinput48 mgmt_gpio_in[20] input48/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XFILLER_155_387 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_115_229 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_109_771 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_124_730 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_96_179 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_4010_ _7720_/Q hold90/I _6107_/A1 _7696_/Q _7680_/Q _6073_/A1 _4013_/A2 VDD VSS
+ gf180mcu_fd_sc_mcu7t5v0__aoi222_1
XFILLER_38_747 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_18_471 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5961_ _7623_/Q _5970_/A2 _5962_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_4912_ _4922_/A3 _4922_/A4 _4924_/A1 _4924_/A2 _4914_/A4 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand4_2
X_7700_ _7700_/D _7923_/RN _7791_/CLK _7700_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffsnq_1
XFILLER_52_238 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_7631_ hold73/Z _7853_/RN _7747_/CLK _7631_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
X_5892_ _4460_/Z _5902_/A2 _5892_/B hold426/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_61_772 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_61_783 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_4843_ _4843_/A1 _6537_/A2 _4847_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_33_496 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_147_800 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_7562_ _7562_/D _7900_/RN _7881_/CLK _7562_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
X_4774_ _4774_/A1 _6537_/A2 _4778_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_3725_ _5006_/C _5254_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__inv_8
XFILLER_158_181 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_146_321 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6513_ _6547_/A1 _6519_/A2 _6513_/B hold443/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_20_179 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_7493_ _7493_/D _7503_/CLK _7493_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_6444_ hold59/Z _6451_/A2 hold60/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_107_708 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3656_ _7915_/Q _6905_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_2
XFILLER_161_357 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6375_ hold64/Z _6383_/A2 _6375_/B _7817_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_5326_ _5326_/A1 _5326_/A2 _5326_/A3 _5326_/A4 _5354_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand4_1
XFILLER_0_529 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_142_593 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_130_744 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5257_ _5394_/A1 _5005_/Z _5622_/A1 _5721_/C VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor3_1
XFILLER_130_788 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_102_479 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4208_ hold942/Z _4427_/B _4284_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_5188_ _5739_/A1 _5188_/A2 _5188_/A3 _5188_/A4 _5191_/B2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand4_1
XFILLER_68_371 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4139_ hold82/Z _4151_/A2 _4599_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_56_566 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_28_268 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_37_780 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_43_227 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_24_463 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_7829_ _7829_/D _7877_/RN _7829_/CLK _7829_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_51_282 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_165_641 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_164_140 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_137_354 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_22_53 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_180_622 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_118_2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_105_240 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_79_636 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_78_124 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_94_617 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_93_105 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_78_179 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_74_330 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_35_706 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_62_514 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_34_205 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_74_396 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1150 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1183 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1172 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1161 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_15_496 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_43_783 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_147_107 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1194 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_8_33 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_128_321 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
Xhold607 _7343_/Q hold607/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
XFILLER_156_685 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xhold618 _7459_/Q hold618/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
X_4490_ _6539_/A1 _4504_/A2 _4490_/B hold843/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
Xmax_cap348 hold63/Z hold64/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__buf_12
XFILLER_143_357 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
Xhold629 hold629/I _7694_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
XFILLER_116_549 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
Xmax_cap359 input75/Z _7961_/RN VDD VSS gf180mcu_fd_sc_mcu7t5v0__buf_20
XFILLER_170_176 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6160_ hold47/Z _6174_/A2 _6160_/B _7716_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
XTAP_901 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_5111_ _5797_/B _5797_/C _5793_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_4
XFILLER_124_593 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_112_744 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_33_2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_912 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_923 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_934 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_6091_ hold620/Z _6106_/A2 hold621/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_945 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_956 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_967 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_978 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_5042_ _5548_/A1 _5043_/A2 _5042_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_97_499 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_84_105 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_989 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_93_650 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_38_544 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_38_566 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_53_503 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xclkbuf_leaf_51_csclk clkbuf_3_6__f_csclk/Z _7818_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
X_6993_ _7831_/Q _7203_/A2 _7204_/B1 _7767_/Q _6997_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_5944_ hold251/Z _5953_/A2 _5945_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_41_709 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_178_210 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5875_ hold487/Z _5880_/A2 _5876_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_80_388 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_21_411 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_21_422 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_7614_ _7614_/D _7923_/RN _7737_/CLK _7614_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
X_4826_ _4826_/A1 _4828_/S _4826_/B _7500_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_7545_ _7545_/D _7959_/RN _7545_/CLK hold52/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
Xclkbuf_leaf_66_csclk clkbuf_3_3__f_csclk/Z _7606_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_147_641 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_119_354 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_21_499 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4757_ hold853/Z _4758_/A2 _4758_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_174_460 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_162_611 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_146_162 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_4688_ _3819_/Z hold47/Z _4689_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_7476_ _7476_/D _7938_/RN _7531_/CLK _7476_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
X_3708_ _7639_/Q _3708_/ZN VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_3639_ _7414_/Q _4383_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_3
X_6427_ hold448/Z _6434_/A2 _6428_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_6358_ hold64/Z _6366_/A2 _6358_/B hold83/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_134_368 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5309_ _5309_/A1 _3723_/I _5344_/A1 _5422_/B _5495_/B2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand4_4
XFILLER_130_530 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6289_ hold168/Z _6298_/A2 _6290_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_88_455 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_88_444 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_124_33 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_102_265 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_84_37 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_90_108 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_84_59 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_72_812 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_56_374 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
Xclkbuf_leaf_19_csclk _7873_/CLK _7899_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_56_396 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_56_385 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_200 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_25_761 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_233 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_222 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_211 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_25_783 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_277 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_266 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_255 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_244 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_157_438 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_299 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_288 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_12_477 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_153_622 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_137_173 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_153_633 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_152_121 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_180_463 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_165_73 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_152_154 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_125_357 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_4_676 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xhold4 hold4/I hold4/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
XFILLER_94_425 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_79_499 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_66_116 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_66_105 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_58_60 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_75_672 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_63_812 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3990_ _3990_/A1 _3990_/A2 _3990_/A3 _3999_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor3_2
XFILLER_62_388 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5660_ _5079_/Z _5660_/A2 _5485_/B _5661_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor3_1
XFILLER_176_747 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4611_ _6539_/A1 _4613_/A2 _4611_/B _7407_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_175_246 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5591_ _5474_/B _5591_/A2 _5454_/B _5656_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor3_1
XFILLER_129_641 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7330_ _7901_/RN _4334_/Z _7330_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__and2_1
X_4542_ hold16/Z _4548_/A2 _4542_/B hold56/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_156_460 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_129_696 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7261_ _7261_/A1 _7261_/A2 _7262_/C VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_143_121 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_116_346 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
Xhold426 hold426/I _7590_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
Xhold415 _8006_/I hold415/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
X_4473_ hold733/Z _4487_/A1 _4477_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
Xhold404 hold404/I _7525_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
Xhold459 hold459/I _6494_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
XFILLER_89_219 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
Xhold448 _7842_/Q hold448/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
Xhold437 _7770_/Q hold437/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
X_6212_ hold928/Z _6225_/A2 _6213_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_171_496 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7192_ _7192_/A1 _7192_/A2 _7192_/A3 _7209_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand3_1
X_6143_ hold47/Z _6157_/A2 _6143_/B hold496/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
XTAP_720 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_731 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_742 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_85_425 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6074_ hold363/Z _6089_/A2 hold364/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_753 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_764 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_775 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_786 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_5025_ _5369_/B _5024_/Z _5535_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_100_747 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_797 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_72_119 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_72_108 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_54_812 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1919 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1908 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_6976_ _6976_/A1 _6976_/A2 _6976_/A3 _6976_/A4 _6977_/A4 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand4_1
X_5927_ hold152/Z _5936_/A2 hold153/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_70_17 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_139_449 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5858_ _6547_/A1 _5868_/A2 _5858_/B _7575_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_5789_ _5789_/A1 _5789_/A2 _5790_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_4809_ _7228_/I0 _7492_/Q _4809_/S _7492_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_135_611 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_119_44 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7528_ _7528_/D _7938_/RN _7528_/CLK _7528_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_147_493 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_7459_ _7459_/D _7853_/RN _7818_/CLK _7459_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_119_55 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_162_463 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_107_357 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xhold960 _7971_/Q hold960/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
XFILLER_134_176 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_89_753 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_89_764 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_123 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_76_425 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_48_105 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_88_296 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_91_428 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_28_52 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_29_363 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_45_812 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_71_141 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_60_804 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_17_558 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_158_703 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_13_753 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_158_747 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_12_263 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_8_201 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_173_706 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_158_758 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_138_460 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_9_779 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_8_256 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_181_783 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_125_132 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_4_451 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_180_282 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_153_496 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_125_176 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_4_473 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_69_70 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_140_179 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_95_712 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_79_296 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_690 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_85_80 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_67_469 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_36_812 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_54_108 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_75_480 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_35_300 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6830_ _7739_/Q _6878_/A2 _6830_/B _6834_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_6761_ _7802_/Q _6883_/A2 _6883_/B1 _7786_/Q _6763_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_3973_ _7380_/Q hold55/I _6282_/A1 _7779_/Q _3985_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_5712_ _5104_/B _5669_/B _5712_/B _5716_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_50_325 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6692_ _6692_/A1 _6692_/A2 _6692_/A3 _6692_/A4 _6706_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand4_1
X_5643_ _5669_/B _5643_/A2 _5643_/B1 _5690_/A1 _5644_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_157_780 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5574_ _5705_/A2 _4996_/Z _5624_/A1 _5624_/B _5736_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_163_238 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xhold201 hold201/I _7699_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
X_4525_ hold856/Z _4526_/A2 _4526_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_7313_ _7900_/RN _4334_/Z _7313_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__and2_1
Xhold234 hold234/I _7754_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
Xhold223 hold223/I _6153_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
XFILLER_144_463 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
Xhold212 hold212/I _7707_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
X_7244_ _7518_/Q _7244_/A2 _7246_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_171_282 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_116_176 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xhold245 _7789_/Q hold245/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
Xhold256 hold256/I _6536_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
Xhold267 hold267/I _7885_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
Xhold278 hold278/I _6534_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
X_4456_ _4487_/A1 _4454_/Z _4456_/B _7348_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_131_146 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4387_ _7448_/Q input89/Z _4387_/S _4387_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
Xhold289 hold289/I _6398_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
X_7175_ _7476_/Q _7195_/A2 _7195_/B1 _7470_/Q _7195_/C1 _7383_/Q _7177_/A3 VDD VSS
+ gf180mcu_fd_sc_mcu7t5v0__aoi222_1
XTAP_550 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_561 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_6126_ hold47/Z _6140_/A2 _6126_/B hold668/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_100_544 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_572 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_583 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_594 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_105_79 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_100_566 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_100_555 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6057_ hold676/Z _6072_/A2 _6058_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_5008_ _5200_/B _5230_/A1 _5024_/A2 _5011_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor3_1
XFILLER_73_428 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_26_300 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1705 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_81_450 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_1749 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1738 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1727 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1716 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_6959_ _6959_/A1 _6959_/A2 _6959_/A3 _6959_/A4 _6977_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand4_1
XFILLER_179_382 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_139_246 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_10_734 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_155_728 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_5_237 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_5_215 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_163_783 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_135_496 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_123_625 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_100_2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_122_124 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xhold790 _7758_/Q hold790/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
XFILLER_122_179 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_77_712 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_162_52 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_76_233 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_39_73 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_77_778 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_18_812 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_36_108 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_17_311 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_29_171 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_72_450 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_45_664 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_60_601 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_44_174 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_177_308 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_60_634 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_32_336 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
Xclkbuf_2_0__f_mgmt_gpio_in[4] clkbuf_0_mgmt_gpio_in[4]/Z _4418_/I1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_71_82 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_158_577 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_146_739 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_146_717 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_161_709 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_126_463 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
Xoutput306 _4424_/Z spimemio_flash_io0_di VDD VSS gf180mcu_fd_sc_mcu7t5v0__buf_4
Xoutput317 _7493_/Q wb_dat_o[15] VDD VSS gf180mcu_fd_sc_mcu7t5v0__buf_4
X_4310_ _7339_/Q _4294_/Z _4311_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_5290_ _5687_/C _5350_/A3 _5290_/B _5291_/C VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi21_1
Xoutput328 _7943_/Q wb_dat_o[25] VDD VSS gf180mcu_fd_sc_mcu7t5v0__buf_4
Xoutput339 _7502_/Q wb_dat_o[6] VDD VSS gf180mcu_fd_sc_mcu7t5v0__buf_4
XFILLER_87_509 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_4241_ _7806_/Q _6350_/A1 _6124_/A1 _7700_/Q _4243_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_141_499 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_113_168 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_68_756 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4172_ _7717_/Q hold90/I _4863_/A1 _7526_/Q _4174_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_67_266 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_55_406 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_36_620 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7931_ _7931_/D _7938_/RN _7938_/CLK _7931_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_55_428 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_82_247 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_24_804 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_36_631 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_35_141 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_35_152 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7862_ _7862_/D _7900_/RN _7862_/CLK _7862_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffsnq_1
X_7793_ _7793_/D _7877_/RN _7829_/CLK _7793_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
X_6813_ _7381_/Q _6882_/A2 _6894_/C1 _7836_/Q _6813_/C _6815_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi221_1
X_6744_ _7841_/Q _6894_/A2 _6659_/Z _7623_/Q _6747_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_3956_ _4206_/A1 _7228_/I0 _3958_/B1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_149_555 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_6675_ _7692_/Q _6881_/B1 _6882_/B1 _7652_/Q _6885_/B1 _7708_/Q _6677_/A3 VDD VSS
+ gf180mcu_fd_sc_mcu7t5v0__aoi222_1
XFILLER_136_205 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_5626_ _5391_/B _5706_/A2 _5626_/A3 _5625_/Z _5726_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand4_1
X_3887_ hold609/Z _3847_/Z _6537_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_4
X_5557_ _5557_/A1 _5557_/A2 _5557_/A3 _5557_/A4 _5557_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__or4_1
XFILLER_117_463 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_3_708 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_151_219 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_145_783 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_117_496 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_117_474 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5488_ _5648_/A1 _5669_/B _5431_/B _5648_/B2 _5803_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_4508_ hold907/Z _4521_/A2 hold908/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_4439_ _7519_/Q _4338_/Z _7513_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_160_764 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_160_742 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7227_ _7227_/I0 _7947_/Q _7228_/S _7947_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_120_617 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_116_34 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_104_179 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_59_712 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7158_ _7158_/A1 _7158_/A2 _7158_/A3 _7158_/A4 _7159_/A4 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand4_1
XFILLER_86_531 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_112_190 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_7089_ _7089_/A1 _7089_/A2 _7089_/A3 _7089_/A4 _7106_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand4_1
XFILLER_100_330 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_59_778 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_391 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_380 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_6109_ hold47/Z _6123_/A2 _6109_/B hold681/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_100_396 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_18_108 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_58_277 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2225 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2214 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2203 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2269 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2258 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2247 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2236 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1524 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1513 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1502 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_92_37 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XPHY_20 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_31 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_1557 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1546 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1535 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_81_280 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_14_314 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_42 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_25_31 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_26_185 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_53 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_64 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_148_2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1579 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1568 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_75 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_41_144 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_86 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_97 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_22_380 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_10_531 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_155_547 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_127_227 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_10_586 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_182_366 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_108_452 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_182_399 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_108_463 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_110_105 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_173_73 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_123_499 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_110_116 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_92_534 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_37_428 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_49_277 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_92_567 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_17_141 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_45_461 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3810_ hold80/Z _3808_/Z _3810_/S hold81/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_21_807 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4790_ _7223_/A1 _4795_/S _4790_/B _7480_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_3741_ _3734_/Z _3741_/A2 _3741_/B _7978_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_60_497 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_174_812 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3672_ _3672_/I _7268_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_6460_ _6545_/A1 _6468_/A2 _6460_/B hold162/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_173_366 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6391_ hold461/Z _6400_/A2 hold462/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_5411_ _5669_/A1 _5793_/A2 _5292_/B _5482_/B2 _5411_/C _5413_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi221_1
XFILLER_63_2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_127_783 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_126_260 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5342_ _5621_/B _5724_/A2 _5759_/C _5721_/B _5343_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XFILLER_99_144 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_142_764 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5273_ _5273_/A1 _5350_/A3 _5793_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_7012_ _7888_/Q _7196_/A2 _7196_/B1 _7638_/Q _7014_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_1
Xoutput169 _4432_/Z irq[1] VDD VSS gf180mcu_fd_sc_mcu7t5v0__buf_4
XFILLER_101_138 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_99_199 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_68_531 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4224_ _7854_/Q _6452_/A1 _6333_/A1 _7798_/Q _4264_/A4 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_4155_ hold609/Z _4155_/A2 _4527_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_110_672 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_95_361 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_56_726 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4086_ _7622_/Q _5954_/A1 _4231_/B1 input58/Z _4092_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_83_567 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_83_589 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7914_ _7914_/D _7923_/RN _7935_/CLK _7914_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_4
XFILLER_70_206 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_36_450 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7845_ _7845_/D _7901_/RN _7864_/CLK _7845_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_168_105 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_23_144 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_149_330 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7776_ _7776_/D _7877_/RN _7877_/CLK _7776_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffsnq_1
X_4988_ _5104_/B _5735_/A2 _5669_/A1 _5705_/A2 _4999_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_149_352 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6727_ _7800_/Q _6883_/A2 _6893_/B1 _7768_/Q _6891_/A2 _7824_/Q _6728_/A4 VDD VSS
+ gf180mcu_fd_sc_mcu7t5v0__aoi222_1
X_3939_ _7812_/Q _6350_/A1 _5971_/A1 _7634_/Q _3940_/A4 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_137_525 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6658_ _6878_/A2 _6658_/A2 _6658_/A3 _6892_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor3_4
XFILLER_125_709 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5609_ _5657_/A4 _5799_/A2 _5609_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_11_33 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_133_720 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6589_ _6590_/A1 _6665_/A2 _6830_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__and2_2
XFILLER_133_731 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_87_26 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_105_499 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_120_469 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_143_65 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_86_383 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_86_372 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_19_428 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2000 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_74_534 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_46_247 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2022 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2033 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2011 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_61_217 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2077 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2066 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2055 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2044 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1332 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1321 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1310 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_27_494 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2099 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2088 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1365 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1354 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1343 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1398 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1387 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1376 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_14_188 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_174_108 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_168_650 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_156_812 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_7_800 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_30_648 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
Xinput27 mask_rev_in[30] input27/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyb_1
Xinput16 mask_rev_in[20] input16/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XFILLER_155_366 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xinput38 mgmt_gpio_in[11] input38/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyb_1
Xinput49 mgmt_gpio_in[21] input49/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XFILLER_6_321 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_182_174 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_109_783 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_170_347 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_136_591 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_124_742 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_151_550 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_124_764 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_111_425 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_2_593 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_35_6 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_96_169 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_77_70 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_77_81 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_65_523 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_37_247 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_80_515 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_65_567 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5960_ _4460_/Z _5970_/A2 _5960_/B _7622_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_4911_ _4924_/A3 _4924_/A4 _3727_/I _4914_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand3_2
X_5891_ hold424/Z _5902_/A2 hold425/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_7630_ _7630_/D _7877_/RN _7752_/CLK _7630_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffsnq_2
X_4842_ _4376_/B _5520_/C _7279_/A2 _4842_/A4 _7506_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand4_1
XFILLER_60_250 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_159_661 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_147_812 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4773_ _4454_/Z _4773_/A2 _4773_/B _7473_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_7561_ _7561_/D _7875_/RN _7563_/CLK _7561_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
X_3724_ _5006_/B _5394_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__inv_3
X_6512_ hold441/Z _6519_/A2 hold442/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_7492_ _7492_/D _7503_/CLK _7492_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_173_141 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6443_ _6545_/A1 _6451_/A2 _6443_/B _7849_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_3655_ _7914_/Q _6908_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__inv_2
X_6374_ hold101/Z _6383_/A2 _6375_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_130_701 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5325_ _5624_/B _5624_/A2 _5724_/A2 _5685_/B _5326_/A4 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_5256_ _5714_/B1 _5622_/A1 _5731_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_102_425 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_102_469 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4207_ _4207_/I0 hold948/Z _4427_/B _7549_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_5187_ _5187_/A1 _5499_/A1 _5187_/A3 _5187_/A4 _5188_/A4 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor4_1
XFILLER_28_236 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_28_247 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4138_ _7741_/Q hold43/I _4559_/A1 _7388_/Q _4158_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_56_534 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4069_ _4069_/A1 _4069_/A2 _7224_/I0 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_2
XFILLER_169_425 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7828_ _7828_/D _7901_/RN _7866_/CLK _7828_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_24_475 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_156_108 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_138_812 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7759_ _7759_/D _7875_/RN _7862_/CLK _7759_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffsnq_1
XFILLER_22_32 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_138_76 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_98_58 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_121_712 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_121_701 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_3_357 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_120_211 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_120_266 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_93_139 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_47_73 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_47_567 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_28_792 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1140 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1173 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1162 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1151 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_15_486 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_42_250 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_129_812 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1195 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1184 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_175_428 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_155_141 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_7_641 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xhold608 _3812_/Z hold608/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
Xmax_cap349 hold47/Z _6539_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__buf_16
Xhold619 hold619/I _7425_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
XFILLER_109_580 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_97_401 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6090_ _6090_/A1 _7285_/A2 _6106_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_4
XFILLER_88_91 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5110_ _4996_/Z _5672_/A2 _5586_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_902 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_913 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_924 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_935 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_5041_ _5024_/Z _5041_/A2 _5533_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_112_767 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_946 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_957 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_968 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_26_2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_979 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_38_534 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xclkbuf_0_wb_clk_i wb_clk_i clkbuf_0_wb_clk_i/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_80_301 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_65_353 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_65_342 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_53_515 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_92_183 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6992_ _6992_/A1 _6992_/A2 _6992_/A3 _6992_/A4 _7001_/B1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand4_1
XFILLER_179_712 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5943_ _4460_/Z _5953_/A2 _5943_/B _7614_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_5874_ _5874_/A1 _7285_/A2 _5880_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_2
XFILLER_61_570 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_138_108 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4825_ _7500_/Q _4828_/S _4826_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_21_434 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_33_283 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7613_ _7613_/D _7938_/RN _7639_/CLK _7613_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_178_277 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_7544_ _7544_/D _7959_/RN _7545_/CLK hold36/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
X_4756_ _6539_/A1 _4758_/A2 _4756_/B _7466_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_4687_ hold560/Z _4718_/A1 hold561/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_3707_ hold78/I _3707_/ZN VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_7475_ _7475_/D _7875_/RN _7822_/CLK _7475_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
X_3638_ hold49/Z _3810_/S VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_12
X_6426_ _6545_/A1 _6434_/A2 _6426_/B _7841_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_162_689 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_161_144 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6357_ _7809_/Q _6366_/A2 _6358_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_161_177 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5308_ _5498_/A2 _5687_/B _5510_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_103_712 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6288_ _4460_/Z _6298_/A2 _6288_/B _7776_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_349 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_130_575 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5239_ _5563_/B2 _5622_/A1 _5572_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_68_191 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_29_534 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_84_673 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_83_150 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_29_567 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_140_33 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_201 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_234 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_223 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_212 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_24_250 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XPHY_267 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_256 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_245 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_157_428 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_289 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_278 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_130_2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_12_456 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_149_86 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_137_130 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_180_420 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_152_166 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_3_154 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_165_85 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_181_73 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xhold5 hold5/I hold5/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
XFILLER_90_632 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_62_323 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_90_676 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_16_784 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_43_570 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_15_283 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_30_242 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4610_ hold914/Z _4613_/A2 _4611_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_5590_ _5582_/Z _5590_/A2 _5590_/B _5639_/C VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_4541_ _7379_/Q _4548_/A2 _4542_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_156_450 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7260_ _7520_/Q _7260_/A2 _7260_/B1 _7519_/Q _7261_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_1
Xhold427 _7858_/Q hold427/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
Xhold405 _7533_/Q hold405/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
X_4472_ _4487_/A1 _6547_/A1 _4472_/B _7351_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
Xhold416 hold416/I _4725_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
XFILLER_143_144 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6211_ _6539_/A1 _6225_/A2 _6211_/B _7740_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
Xhold449 _7826_/Q hold449/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
Xhold438 _7890_/Q hold438/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
X_7191_ _7510_/Q _7191_/A2 _7191_/B1 _7406_/Q _7192_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_143_177 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6142_ hold494/Z _6157_/A2 hold495/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_112_520 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_98_732 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_710 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_112_531 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_721 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_732 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_743 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_112_564 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6073_ _6073_/A1 _7285_/A2 _6089_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_4
XFILLER_97_286 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_754 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_765 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_776 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_5024_ _3728_/I _5024_/A2 _5024_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__xor2_1
XTAP_798 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_787 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_66_673 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_53_323 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1909 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_53_345 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6975_ _7830_/Q _7203_/A2 _7204_/A2 _7838_/Q _6976_/A4 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_5926_ _4460_/Z _5936_/A2 _5926_/B _7606_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_110_47 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_139_439 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_139_428 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5857_ hold385/Z _5868_/A2 _5858_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_166_247 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5788_ _5412_/B _5788_/A2 _5789_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_21_286 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_4808_ _7227_/I0 _7491_/Q _4809_/S _7491_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_166_269 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4739_ hold730/Z _4750_/I1 _4741_/S _7455_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_119_141 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_119_23 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7527_ _7527_/D _7938_/RN _7961_/CLK _7527_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
X_7458_ _7458_/D _7853_/RN _7601_/CLK _7458_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
X_6409_ _6545_/A1 _6417_/A2 _6409_/B _7833_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
Xhold961 _3767_/Z _7971_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
Xhold950 _7343_/Q hold950/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
XFILLER_134_188 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7389_ _7389_/D _7875_/RN _7637_/CLK _7389_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_135_33 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_115_380 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_103_531 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_103_520 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_135_88 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_135_66 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_89_798 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_95_59 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_28_64 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_29_353 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_178_2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_57_695 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_44_356 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_72_676 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_25_570 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_44_389 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_157_247 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_13_798 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_40_595 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_172_206 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_60_51 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_60_62 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_180_250 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_125_144 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_5_24 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xclkbuf_leaf_50_csclk clkbuf_3_7__f_csclk/Z _7600_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_4_463 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_140_125 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_95_702 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_95_757 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_94_212 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_79_286 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_39_139 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
Xclkbuf_leaf_65_csclk clkbuf_3_3__f_csclk/Z _7791_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_85_70 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_85_92 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_48_673 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_47_194 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_90_473 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_6760_ _7842_/Q _6894_/A2 _6891_/A2 _7826_/Q _6763_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_62_175 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5711_ _5711_/A1 _5733_/A3 _5710_/Z _5717_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand3_1
X_3972_ _7360_/Q _4488_/A1 _6401_/A1 _7835_/Q _3996_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_93_2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_90_495 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6691_ _7759_/Q _6892_/A2 _6893_/C1 _7629_/Q _6692_/A4 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_176_534 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_148_247 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5642_ _5642_/A1 _5642_/A2 _5642_/A3 _5642_/A4 _5766_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand4_1
XFILLER_176_578 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5573_ _5573_/A1 _5759_/A1 _5573_/B _5573_/C _5732_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XFILLER_156_280 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xhold202 _7805_/Q hold202/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
X_4524_ _6539_/A1 _4526_/A2 _4524_/B _7371_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_7312_ _7900_/RN _4334_/Z _7312_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__and2_1
Xhold224 hold224/I _7713_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
Xhold235 _7811_/Q hold235/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
Xhold213 _7739_/Q hold213/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
X_7243_ _7243_/A1 _7277_/B _7243_/B _7950_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_171_272 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4455_ _4455_/A1 hold12/Z hold13/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
Xhold246 _7837_/Q hold246/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
Xhold268 _7901_/Q hold268/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
Xhold257 hold257/I _7893_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
X_4386_ _7449_/Q input91/Z _4387_/S _4386_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_7174_ _7523_/Q _7194_/A2 _7194_/B1 _7504_/Q _7194_/C1 _7409_/Q _7177_/A2 VDD VSS
+ gf180mcu_fd_sc_mcu7t5v0__aoi222_1
Xhold279 hold279/I _7892_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
XTAP_540 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_551 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_6125_ hold666/Z _6140_/A2 hold667/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_112_394 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_100_534 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_85_212 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_562 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_573 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_584 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_595 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_27_802 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6056_ _6056_/A1 _7285_/A2 _6072_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_4
X_5007_ _4898_/Z _4915_/Z _5005_/Z _5151_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand3_2
XFILLER_54_621 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1706 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1739 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1728 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1717 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_121_68 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_81_473 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_81_462 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_54_676 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_81_495 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6958_ _7774_/Q _7200_/A2 _7189_/B1 _7684_/Q _7195_/B1 _7620_/Q _6959_/A4 VDD VSS
+ gf180mcu_fd_sc_mcu7t5v0__aoi222_1
XFILLER_41_337 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_41_348 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5909_ _4460_/Z _5919_/A2 _5909_/B hold493/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_6889_ _7526_/Q _6889_/A2 _6665_/Z _7538_/Q _6889_/C _6896_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi221_1
XFILLER_167_556 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_22_584 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_22_595 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_148_770 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_182_559 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_108_623 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_107_144 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_162_250 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_150_401 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_123_637 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
Xhold791 _7534_/Q hold791/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
Xhold780 _7391_/Q hold780/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
XFILLER_103_361 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_1_499 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_39_52 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_76_245 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_92_738 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_91_215 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_29_150 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_57_481 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_72_473 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_60_613 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_55_73 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_158_534 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_40_392 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_139_792 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
Xoutput307 _4425_/ZN spimemio_flash_io1_di VDD VSS gf180mcu_fd_sc_mcu7t5v0__buf_4
XFILLER_181_570 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_114_626 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_114_615 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
Xoutput329 _7944_/Q wb_dat_o[26] VDD VSS gf180mcu_fd_sc_mcu7t5v0__buf_4
XFILLER_5_783 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_5_772 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
Xoutput318 _7478_/Q wb_dat_o[16] VDD VSS gf180mcu_fd_sc_mcu7t5v0__buf_4
XFILLER_153_283 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4240_ _4240_/A1 _4240_/A2 _4240_/A3 _4240_/A4 _4283_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand4_2
X_4171_ _7522_/Q _4853_/A1 _4873_/A1 _7530_/Q _4174_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_67_212 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_95_576 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7930_ _7930_/D _7961_/RN _7940_/CLK _7930_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
X_7861_ _7861_/D _7901_/RN _7869_/CLK _7861_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
X_6812_ _6812_/A1 _6812_/A2 _6812_/A3 _6813_/C VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_36_676 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_51_602 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7792_ _7792_/D _7923_/RN _7792_/CLK _7792_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffsnq_1
XFILLER_23_337 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_149_512 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6743_ _7615_/Q _6647_/Z _6887_/B1 _7679_/Q _6752_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_3955_ _3955_/A1 _3955_/A2 _3936_/Z _3955_/A4 _7228_/I0 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand4_4
XFILLER_51_668 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6674_ _7782_/Q _6883_/B1 _6891_/C1 _7774_/Q _6674_/C _6677_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi221_1
XFILLER_176_353 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_164_504 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_149_567 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3886_ hold38/Z _3886_/A2 _5988_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_4
X_5625_ _5803_/A2 _5625_/A2 _5625_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__and2_1
X_5556_ _5642_/A4 _5649_/A4 _5557_/A4 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_144_250 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5487_ _5099_/B _5797_/A2 _5645_/A3 _5495_/B2 _5511_/C VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai22_1
X_4507_ _6539_/A1 _4521_/A2 _4507_/B hold849/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_172_592 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4438_ _5678_/A1 _4438_/A2 _7514_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_7226_ _7226_/A1 _7228_/S _7226_/B _7946_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_120_607 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4369_ input97/Z input96/Z input99/Z input98/Z _4374_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor4_1
X_7157_ _7765_/Q _7202_/C2 _7200_/B1 _7869_/Q _7158_/A4 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_98_392 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7088_ _7713_/Q _7189_/A2 _7191_/B1 _7803_/Q _7089_/A4 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XTAP_392 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_370 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_381 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_6108_ hold679/Z _6123_/A2 hold680/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_132_34 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6039_ _6039_/A1 hold5/Z _6055_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_4
XFILLER_73_215 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_46_429 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2226 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2215 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2204 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2259 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2248 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2237 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1514 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1503 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_21 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_10 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_42_602 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1547 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1536 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1525 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_81_292 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_81_270 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_32 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_43 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_54 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_65 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_41_101 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1569 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1558 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_76 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_87 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_98 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_167_375 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_10_521 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_22_392 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_6_514 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_41_75 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_182_356 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_108_431 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_163_570 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_135_294 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_135_283 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_151_776 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_96_318 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_1_241 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_96_329 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_49_212 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_1_296 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_2_47 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_49_256 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_92_546 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_18_676 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_72_270 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_159_810 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_60_443 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_3740_ _4292_/B _3738_/Z _3741_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_60_487 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3671_ _3671_/I _7263_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_118_206 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_9_374 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5410_ _5669_/A1 _5793_/A2 _5292_/B _5482_/B2 _5794_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_6390_ _4460_/Z _6400_/A2 _6390_/B _7824_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_126_250 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_114_412 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5341_ _5645_/A3 _5495_/B2 _5721_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_56_2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_142_754 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_5_580 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5272_ _5199_/B _5201_/B _5338_/A1 _5369_/B _5350_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand4_4
X_7011_ _7646_/Q _7195_/A2 _7195_/B1 _7622_/Q _7188_/A2 _7377_/Q _7016_/A3 VDD VSS
+ gf180mcu_fd_sc_mcu7t5v0__aoi222_1
XFILLER_141_286 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4223_ _7838_/Q _6418_/A1 _4579_/A1 _7395_/Q _4256_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_4154_ hold609/Z _3881_/Z _5807_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_4085_ _7686_/Q _6090_/A1 hold150/I _7565_/Q _6141_/A1 _7710_/Q _4092_/A2 VDD VSS
+ gf180mcu_fd_sc_mcu7t5v0__aoi222_2
XFILLER_28_407 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_55_215 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_7913_ _7913_/D _7923_/RN _7935_/CLK _7913_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_4
XFILLER_102_37 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_24_602 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7844_ _7844_/D _7901_/RN _7858_/CLK _7844_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_24_646 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_51_410 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_169_618 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_23_123 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_24_657 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7775_ _7775_/D _7875_/RN _7863_/CLK _7775_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffsnq_1
X_4987_ _5669_/A1 _5705_/A2 _5706_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_6726_ _7792_/Q _6893_/A2 _6892_/B1 _7726_/Q _6890_/B1 _7848_/Q _6728_/A3 VDD VSS
+ gf180mcu_fd_sc_mcu7t5v0__aoi222_1
XFILLER_51_487 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_165_802 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3938_ input41/Z _5903_/A1 _6039_/A1 _7666_/Q _3940_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_3869_ _3869_/I _4653_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_6657_ _6878_/A2 _6661_/A3 _6658_/A3 _6893_/B1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor3_4
XFILLER_176_194 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5608_ _5608_/A1 _5167_/B _5608_/B _5799_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_6588_ _7909_/Q _7908_/Q _6665_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_2
XFILLER_164_389 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5539_ _5543_/B _5153_/C _5539_/A3 _5552_/A4 _5546_/C VDD VSS gf180mcu_fd_sc_mcu7t5v0__or4_1
XFILLER_152_529 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_145_570 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_117_283 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_87_16 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_79_808 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_11_89 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_78_318 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_143_11 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_132_275 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_59_510 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7209_ _7210_/A2 _7209_/A2 _7209_/A3 _7209_/A4 _7210_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor4_1
XFILLER_59_554 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_100_150 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_74_513 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_46_204 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2001 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_100_183 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2023 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2034 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2012 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_160_2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2067 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2056 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2045 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1322 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1311 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1300 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2089 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2078 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1366 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1355 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1344 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1333 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_14_134 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_30_605 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1399 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1388 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1377 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_52_41 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_168_673 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_52_63 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_167_172 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_10_362 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_7_812 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xinput28 mask_rev_in[31] input28/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyb_1
Xinput17 mask_rev_in[21] input17/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XFILLER_182_142 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xinput39 mgmt_gpio_in[12] input39/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyc_1
XFILLER_108_261 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_108_250 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_124_721 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_123_242 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_123_286 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_97_638 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_69_329 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_96_159 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_93_811 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_37_204 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_37_215 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_92_321 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_46_771 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_46_760 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4910_ input97/Z input96/Z input99/Z input98/Z _4914_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand4_4
XFILLER_93_70 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_80_527 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5890_ _4454_/Z _5902_/A2 _5890_/B _7589_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_4841_ hold49/I _7214_/A1 _4842_/A4 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_178_459 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_21_638 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_33_476 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4772_ hold814/Z _4773_/A2 _4773_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_7560_ _7560_/D _7875_/RN _7563_/CLK _7560_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffsnq_1
X_3723_ _3723_/I _5087_/C VDD VSS gf180mcu_fd_sc_mcu7t5v0__inv_4
XFILLER_9_160 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_6511_ _6545_/A1 _6519_/A2 _6511_/B hold146/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_7491_ _7491_/D _7503_/CLK _7491_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_6442_ hold163/Z _6451_/A2 _6443_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_3654_ _7911_/Q _6599_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_2
XFILLER_174_676 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_146_389 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_127_570 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_115_721 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6373_ _4460_/Z _6383_/A2 _6373_/B _7816_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_5324_ _5624_/B _5624_/A2 _5647_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_88_605 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_115_798 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5255_ _5273_/A1 _5687_/C _5705_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_87_159 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_87_148 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4206_ _4206_/A1 _7221_/A1 _4206_/B _4207_/I0 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_5186_ _5186_/A1 _5186_/A2 _5186_/A3 _5186_/A4 _5187_/A4 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand4_1
XFILLER_84_811 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4137_ hold82/Z _4217_/A2 _4559_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_56_546 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_56_557 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4068_ _4068_/A1 _4068_/A2 _4069_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_83_354 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7827_ _7827_/D _7901_/RN _7829_/CLK _7827_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_169_437 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_12_605 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_51_262 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_7758_ _7758_/D _7875_/RN _7862_/CLK _7758_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffsnq_1
X_7689_ _7689_/D _7923_/RN _7698_/CLK _7689_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
X_6709_ _7922_/Q _7133_/S _6710_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_138_33 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_20_671 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_180_602 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_138_66 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_138_55 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_98_26 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_98_37 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_105_242 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_105_286 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_79_638 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_78_104 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_160_392 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_87_682 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_93_129 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_87_693 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_74_321 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_19_215 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_74_376 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_28_782 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1141 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1130 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1174 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1163 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1152 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_63_73 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_179_73 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1196 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1185 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_11_682 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_156_676 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xhold609 hold609/I hold609/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
XFILLER_128_389 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_116_529 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_7_664 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_170_123 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_109_570 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_143_359 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_124_540 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_124_551 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_111_212 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_88_70 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_903 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_914 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_925 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_5040_ _5151_/A1 _5151_/A2 _5040_/B _5043_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi21_2
XFILLER_111_223 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_69_148 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_936 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_947 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_958 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_969 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_93_641 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_77_170 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_19_2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_93_652 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6991_ _6991_/A1 _6991_/A2 _6992_/A4 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_5942_ hold549/Z _5953_/A2 _5943_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_18_270 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_92_195 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_178_212 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5873_ _6539_/A1 _5873_/A2 _5873_/B _7582_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_178_267 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7612_ _7612_/D _7961_/RN _7639_/CLK _7612_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffsnq_1
X_4824_ _7224_/I0 _7499_/Q _4828_/S _7499_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_147_621 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_119_312 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7543_ _7543_/D _7959_/RN _7545_/CLK hold80/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
X_4755_ hold779/Z _4758_/A2 _4756_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_3706_ _7655_/Q _3706_/ZN VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_162_602 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4686_ _4686_/A1 _5903_/A2 _4686_/B1 _3819_/Z hold22/Z _4718_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi221_4
X_7474_ _7474_/D _7875_/RN _7547_/CLK _7474_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
X_3637_ _7344_/Q _3744_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__inv_1
X_6425_ hold167/Z _6434_/A2 _6426_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_150_808 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6356_ _4460_/Z _6366_/A2 _6356_/B _7808_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_108_69 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5307_ _5307_/A1 _5307_/A2 _5650_/A3 _5433_/C _5307_/B2 _5356_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai32_1
XFILLER_115_595 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_102_212 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_317 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_170_690 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_142_392 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6287_ hold694/Z _6298_/A2 _6288_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_103_768 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_5238_ _5200_/B _3727_/I _5421_/A1 _5422_/B _5622_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand4_4
X_5169_ _5643_/A2 _5672_/A2 _5793_/A2 _5167_/B _5171_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_124_79 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_124_68 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_84_17 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_69_693 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_56_321 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_56_332 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_17_708 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_17_33 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_44_538 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_56_398 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_71_357 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_169_212 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_224 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_213 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_202 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_25_763 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_169_245 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_268 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_257 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_246 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_235 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_12_446 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_40_744 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_279 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_137_120 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_123_2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_138_676 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_141_808 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_106_551 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_3_144 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_140_318 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xhold6 hold6/I hold6/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
XFILLER_47_310 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_75_674 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_75_641 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_47_354 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_15_240 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_175_215 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_175_248 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4540_ _6545_/A1 _4548_/A2 _4540_/B _7378_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_144_602 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_144_646 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
Xhold417 hold417/I _7446_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
XFILLER_7_494 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4471_ hold614/Z _4487_/A1 _4472_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
Xhold406 hold406/I _4885_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
X_6210_ hold860/Z _6225_/A2 _6211_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_116_348 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xhold428 hold428/I _6462_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
Xhold439 hold439/I _6530_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
X_7190_ _7402_/Q _7190_/A2 _7190_/B1 _7469_/Q _7190_/C1 _7526_/Q _7192_/A2 VDD VSS
+ gf180mcu_fd_sc_mcu7t5v0__aoi222_1
X_6141_ _6141_/A1 _7285_/A2 _6157_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_4
XTAP_700 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_124_392 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_98_744 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_711 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_722 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_733 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_6072_ _6553_/A1 _6072_/A2 _6072_/B hold198/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_98_788 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_744 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_755 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_766 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_777 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_39_811 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5023_ _5338_/A1 _5024_/A2 _5040_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_85_449 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_799 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_788 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_38_321 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_93_460 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_26_538 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_38_387 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_53_357 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6974_ _7644_/Q _7195_/A2 _7190_/B1 _7612_/Q _6976_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_80_176 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5925_ hold610/Z _5936_/A2 _5926_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_179_565 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_110_37 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5856_ _5870_/A1 _7285_/A2 _5868_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_4
XFILLER_22_733 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_179_587 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4807_ _4826_/A1 _4809_/S _4807_/B _7490_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_21_232 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_5787_ _5787_/A1 _5787_/A2 _5787_/A3 _7544_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_182_719 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_175_771 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_4738_ hold420/Z _4749_/I1 _4741_/S _4738_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_7526_ _7526_/D _7938_/RN _7741_/CLK _7526_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
X_4669_ _4685_/A1 hold465/Z _4669_/B hold466/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_7457_ _7457_/D _7853_/RN _7601_/CLK _7457_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_150_605 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6408_ hold182/Z _6417_/A2 _6409_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
Xhold940 _7551_/Q hold940/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
Xhold962 hold15/I hold962/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
Xhold951 _7415_/Q _3662_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
XFILLER_122_318 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_115_370 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7388_ _7388_/D input75/Z _7477_/CLK _7388_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
X_6339_ _4460_/Z _6349_/A2 _6339_/B _7800_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_1_637 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_130_362 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_88_254 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_158 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8009_ _8009_/I _8009_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_57_641 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_151_44 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_72_611 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_71_154 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_32_519 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_44_368 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_157_215 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_13_777 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_158_749 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_126_602 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_8_247 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_60_41 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_126_646 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_141_638 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_106_392 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_121_373 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_94_202 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_10_6 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_75_460 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_48_696 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_62_110 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3971_ _7899_/Q _6537_/A1 _4719_/A1 _8009_/I _3998_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_90_463 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_35_357 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5710_ _5710_/A1 _5710_/A2 _5710_/A3 _5710_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__and3_1
XFILLER_62_187 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_149_716 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_149_738 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6690_ _7823_/Q _6891_/A2 _6891_/B1 _7669_/Q _6892_/B1 _7725_/Q _6692_/A3 VDD VSS
+ gf180mcu_fd_sc_mcu7t5v0__aoi222_1
X_5641_ _5641_/A1 _5641_/A2 _5558_/B _5747_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_86_2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5572_ _4996_/Z _5608_/B _5572_/B _5572_/C _5716_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi211_2
X_4523_ hold764/Z _4526_/A2 _4524_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_7311_ _7900_/RN _4334_/Z _7311_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__and2_1
X_7242_ _7242_/A1 _7280_/A2 _7277_/B _7242_/C _7243_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XFILLER_172_763 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_172_741 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xhold225 _7665_/Q hold225/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
Xhold203 hold203/I _7805_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
Xhold214 hold214/I _6208_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
XFILLER_171_262 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4454_ _4455_/A1 hold12/Z _4454_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__and2_4
XFILLER_132_605 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xhold236 hold236/I _7811_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
XFILLER_116_156 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
Xhold258 _7781_/Q hold258/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
XFILLER_104_318 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_104_329 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
Xhold269 hold269/I _6553_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
Xhold247 _7358_/Q hold247/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
X_4385_ _5678_/A1 _4338_/Z _7215_/C _7516_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_171_295 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_131_137 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_7173_ _7395_/Q _7193_/A2 _7193_/B1 _7472_/Q _7193_/C1 _7531_/Q _7177_/A1 VDD VSS
+ gf180mcu_fd_sc_mcu7t5v0__aoi222_1
X_6124_ _6124_/A1 _7285_/A2 _6140_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_4
XTAP_530 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_541 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_552 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_6055_ _6553_/A1 _6055_/A2 _6055_/B hold109/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_86_747 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_563 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_574 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_585 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_5006_ _3722_/I _3723_/I _5006_/B _5006_/C _5024_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai211_4
XFILLER_105_59 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_596 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_39_641 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_66_460 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1729 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1718 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1707 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_53_154 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6957_ _7814_/Q _7207_/A2 _7190_/C1 _7700_/Q _6959_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_81_485 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_139_215 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5908_ hold491/Z _5919_/A2 hold492/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_6888_ _6888_/A1 _6888_/A2 _6888_/A3 _6888_/A4 _6888_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__and4_1
XFILLER_139_248 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5839_ hold704/Z _5840_/A2 _5840_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_108_602 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_10_747 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_182_527 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7509_ _7509_/D _7961_/RN _7572_/CLK _7509_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_163_774 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_135_476 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_122_104 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_107_156 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_146_99 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_146_77 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_107_189 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_1_423 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
Xhold770 _7586_/Q hold770/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
Xhold781 _7385_/Q hold781/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
XFILLER_150_479 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
Xhold792 hold792/I _4887_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
XFILLER_1_456 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_103_384 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_89_585 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_77_736 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_49_416 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_92_717 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_17_313 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_72_463 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_17_357 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_72_496 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_60_636 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_44_176 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_71_73 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_9_567 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_138_270 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_138_281 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
Xoutput308 _8008_/Z spimemio_flash_io2_di VDD VSS gf180mcu_fd_sc_mcu7t5v0__buf_4
XFILLER_153_240 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_126_465 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_114_605 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_113_104 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_4_250 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xoutput319 _7479_/Q wb_dat_o[17] VDD VSS gf180mcu_fd_sc_mcu7t5v0__buf_4
XFILLER_58_6 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_153_295 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_99_338 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4170_ _4167_/Z _4170_/A2 _4170_/A3 _4204_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_68_747 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_68_736 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_96_81 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_95_588 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_48_460 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_48_471 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_75_290 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7860_ _7860_/D _7900_/RN _7878_/CLK _7860_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_91_783 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6811_ _7666_/Q _6885_/A2 _6893_/B1 _7772_/Q _6812_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_90_260 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_63_496 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7791_ _7791_/D _7938_/RN _7791_/CLK _7791_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffsnq_1
XFILLER_177_800 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_6742_ _6742_/A1 _6742_/A2 _6742_/A3 _6753_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand3_1
X_3954_ _3954_/A1 _3954_/A2 _3954_/A3 _3954_/A4 _3955_/A4 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor4_4
XFILLER_176_321 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3885_ _3847_/Z hold82/Z _6401_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_4
XFILLER_50_179 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_6673_ _6673_/A1 _6673_/A2 _6673_/A3 _6674_/C VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand3_1
X_5624_ _5624_/A1 _5624_/A2 _5648_/B2 _5624_/B _5626_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai31_1
XFILLER_164_527 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_129_281 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5555_ _5179_/B _5793_/A2 _5555_/B _5555_/C _5649_/A4 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi211_2
X_5486_ _5543_/B _5504_/B1 _5553_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_104_104 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4506_ hold847/Z _4521_/A2 hold848/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_4437_ _7518_/Q _4338_/Z _7515_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_160_744 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_105_638 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7225_ _7946_/Q _7228_/S _7226_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_7156_ _7805_/Q _7191_/B1 _7188_/A2 _7382_/Q _7158_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_4368_ _4368_/A1 _4368_/A2 _4368_/A3 _4372_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor3_1
XFILLER_113_693 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_113_682 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6107_ _6107_/A1 _7285_/A2 _6123_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_4
X_4299_ _7343_/Q _4383_/A1 _4297_/Z _4300_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand3_1
X_7087_ _7689_/Q _7189_/B1 _7189_/C1 _7657_/Q _7089_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_100_321 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_86_566 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_371 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_393 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_382 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_58_246 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_132_13 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6038_ _6553_/A1 _6038_/A2 _6038_/B hold191/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_27_611 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2216 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2205 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_73_227 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_27_622 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_27_633 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2249 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2238 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2227 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1515 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1504 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_22 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_11 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_54_463 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7989_ _7989_/I _7989_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_1548 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1537 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1526 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_33 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_44 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_27_699 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XPHY_55 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_1559 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_25_77 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_66 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_77 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_88 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_99 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_167_354 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xclkbuf_leaf_64_csclk clkbuf_3_3__f_csclk/Z _7733_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_157_43 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_136_741 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_136_763 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_150_210 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_108_498 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_104_682 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_1_286 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_2_37 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_18_666 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
Xclkbuf_leaf_17_csclk _7873_/CLK _7833_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_73_783 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_45_496 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_32_124 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_158_321 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_32_179 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3670_ _3670_/I _7258_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_146_527 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_9_353 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_173_357 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_142_700 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_127_763 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_5340_ _5689_/A2 _5687_/B _5504_/A3 _5618_/B1 _5498_/A2 _5759_/C VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai32_1
XFILLER_142_744 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5271_ _3728_/I _5022_/B _5271_/A3 _5431_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor3_4
XFILLER_99_124 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_5_570 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_49_2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7010_ _7694_/Q _7194_/A2 _7194_/B1 _7662_/Q _7194_/C1 _7808_/Q _7016_/A2 VDD VSS
+ gf180mcu_fd_sc_mcu7t5v0__aoi222_1
X_4222_ _7774_/Q _6282_/A1 _4584_/A1 _7397_/Q _4264_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_4153_ hold38/Z _3959_/Z _4812_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_4084_ _4084_/A1 _4084_/A2 _4084_/A3 _4084_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__and3_1
XFILLER_83_514 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7912_ _7912_/D _7923_/RN _7935_/CLK _7912_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffsnq_4
XFILLER_49_791 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_71_709 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_64_761 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_36_463 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7843_ _7843_/D _7901_/RN _7869_/CLK _7843_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_91_591 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_91_580 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4986_ _4993_/B _5647_/A2 _5705_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_4
X_7774_ _7774_/D _7875_/RN _7863_/CLK _7774_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffsnq_1
X_6725_ _7808_/Q _6880_/B1 _6665_/Z _7742_/Q _6728_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_3937_ _7780_/Q _6282_/A1 _6248_/A1 _7764_/Q _6401_/A1 _7836_/Q _3940_/A2 VDD VSS
+ gf180mcu_fd_sc_mcu7t5v0__aoi222_2
XFILLER_23_157 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_51_499 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_177_641 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_176_140 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_149_354 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_149_332 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3868_ hold26/Z _3925_/A2 hold75/Z _3963_/A4 _3869_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__or4_4
X_6656_ _6878_/A2 _6664_/A3 _6658_/A3 _6891_/C1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor3_4
X_3799_ _7341_/Q _7414_/Q _7342_/Q _3801_/I1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi21_2
X_5607_ _5648_/A2 _5606_/B _5657_/A4 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_6587_ _6636_/A1 _6587_/A2 _6587_/B _7909_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_5538_ _5538_/A1 _5548_/A1 _5643_/B1 _5150_/Z _5652_/A4 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand4_1
XFILLER_117_240 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_5469_ _5735_/A2 _5643_/A2 _5672_/A2 _4996_/Z _5749_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_7208_ _7208_/A1 _7208_/A2 _7208_/A3 _7208_/A4 _7209_/A4 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand4_1
XFILLER_143_45 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_101_641 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7139_ _7821_/Q _7207_/A2 _7201_/A2 _7755_/Q _7140_/A4 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_86_330 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_100_140 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2024 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2013 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2002 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_27_452 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_36_32 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2068 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2057 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2046 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2035 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1323 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1312 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1301 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_27_496 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_55_783 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2079 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_153_2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1356 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1345 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1334 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_14_124 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1389 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1367 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1378 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_14_179 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_128_516 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xinput18 mask_rev_in[22] input18/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyc_1
XFILLER_171_806 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_155_357 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xinput29 mask_rev_in[3] input29/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XFILLER_136_593 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_124_744 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_6_389 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_117_90 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_111_416 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_96_127 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_96_116 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_96_105 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_35_8 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_65_503 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_65_547 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_53_709 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_18_463 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_4840_ _7517_/D _7513_/Q _7515_/Q _7514_/Q _7279_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor4_2
XFILLER_61_753 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_60_263 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_20_105 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_21_628 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_33_466 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_159_641 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1890 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_4771_ _6539_/A1 _4773_/A2 _4771_/B _7472_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_6510_ hold144/Z _6519_/A2 hold145/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_33_499 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_174_600 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3722_ _3722_/I _5309_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_8
X_7490_ _7490_/D _7949_/CLK _7490_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_6441_ _4460_/Z _6451_/A2 _6441_/B _7848_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_146_346 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3653_ _7434_/Q _4352_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_2
XFILLER_174_666 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_173_165 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_161_316 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_134_519 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_134_508 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6372_ hold626/Z _6383_/A2 _6373_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_173_176 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_127_582 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5323_ _5724_/B _5648_/B2 _5724_/A2 _5624_/B _5326_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_5254_ _5006_/B _5254_/A2 _5254_/A3 _5422_/B _5409_/B2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand4_4
XFILLER_87_105 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5185_ _5666_/A1 _5669_/B _5185_/B _5512_/B _5186_/A4 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XFILLER_130_747 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_68_330 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4205_ _7548_/Q _4206_/A1 _4206_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_110_460 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4136_ hold54/Z _4155_/A2 _6243_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_4067_ _4067_/A1 _4067_/A2 _4067_/A3 _4067_/A4 _4068_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand4_1
XFILLER_36_260 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_37_783 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7826_ _7826_/D _7901_/RN _7854_/CLK _7826_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
X_4969_ _5774_/A1 _5709_/A1 _4969_/B _4969_/C _4999_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai211_1
X_7757_ _7757_/D _7875_/RN _7790_/CLK _7757_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
X_7688_ _7688_/D _7923_/RN _7792_/CLK _7688_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_22_34 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6708_ _7433_/Q _7921_/Q _6708_/B _6710_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_6639_ _6878_/A2 _6663_/A4 _6658_/A3 _6883_/B1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor3_4
XFILLER_153_806 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_137_357 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_164_176 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_98_49 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_121_703 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_106_744 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_121_736 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_154_66 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_105_298 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_101_460 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_86_160 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1120 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1131 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_63_30 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_179_30 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1164 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1153 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1142 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1197 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1186 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1175 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_15_499 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_168_460 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_155_132 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_156_666 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_155_165 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_155_176 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_143_316 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_170_179 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_112_736 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_97_403 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_904 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_915 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_926 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_112_747 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_88_93 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_2_392 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_937 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_948 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_959 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_84_108 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_66_812 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_77_160 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_65_300 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6990_ _6990_/A1 _6990_/A2 _6990_/A3 _6990_/A4 _6991_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand4_1
XFILLER_19_761 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_19_783 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5941_ _4454_/Z _5953_/A2 _5941_/B _7613_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_34_742 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_61_550 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5872_ hold751/Z _5873_/A2 _5873_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_166_408 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_7611_ _7611_/D _7923_/RN _7792_/CLK _7611_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
X_4823_ _7223_/A1 _4828_/S _4823_/B _7498_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_147_611 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7542_ _7542_/D _7959_/RN _7545_/CLK hold24/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_119_302 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4754_ _4754_/A1 _6537_/A2 _4758_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_3705_ hold79/I _3705_/ZN VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_7473_ _7473_/D _7961_/RN _7531_/CLK _7473_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_174_463 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_119_357 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_4685_ _4685_/A1 _4685_/A2 _4685_/B hold231/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_146_176 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6424_ _4460_/Z _6434_/A2 _6424_/B _7840_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_3636_ _3636_/I _4002_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_6355_ hold688/Z _6366_/A2 _6356_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_108_37 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_1_808 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5306_ _5645_/A1 _5421_/B1 _5650_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_115_585 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6286_ _4454_/Z _6298_/A2 _6286_/B _7775_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_103_758 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5237_ _5433_/C _5621_/B _5237_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_111_780 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5168_ _5643_/A2 _5672_/A2 _5673_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_96_491 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_96_480 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5099_ _4993_/C _5663_/A1 _5099_/B _5573_/C VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_83_141 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4119_ hold54/Z _4217_/A2 _4604_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_83_163 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_71_347 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_25_753 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XPHY_225 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_214 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_203 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_52_550 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7809_ hold83/Z _7877_/RN _7809_/CLK _7809_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_169_235 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_258 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_247 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_236 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_33_33 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_269 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_12_469 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_40_756 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_177_290 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_33_99 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_153_614 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_138_666 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_126_806 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_180_400 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_165_496 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_116_2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_4_602 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_4_646 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_152_179 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_79_425 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_160_190 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_79_436 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_58_30 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_66_108 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_48_812 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_58_52 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
Xhold7 hold7/I hold7/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
XFILLER_35_506 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_74_196 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_31_712 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_129_611 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_129_633 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_128_121 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_156_463 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_128_143 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xhold418 _7462_/Q hold418/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
X_4470_ hold16/Z _4749_/I1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_128_176 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xhold407 hold407/I _7533_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
XFILLER_99_92 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_99_70 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xhold429 hold429/I _7858_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
XFILLER_171_499 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_143_168 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6140_ _6553_/A1 _6140_/A2 _6140_/B hold212/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
XTAP_701 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_124_382 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_112_544 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_712 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_31_2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_723 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_734 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_6071_ hold196/Z _6072_/A2 hold197/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_97_277 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_745 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_756 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_767 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_5022_ _5338_/A1 _5024_/A2 _5022_/B _5151_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_2
XFILLER_100_739 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_97_288 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_85_428 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_778 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_789 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_65_141 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6973_ _7708_/Q _7189_/A2 _7193_/B1 _7628_/Q _6938_/I _7854_/Q _6976_/A2 VDD VSS
+ gf180mcu_fd_sc_mcu7t5v0__aoi222_1
X_5924_ _4454_/Z _5936_/A2 _5924_/B _7605_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_41_509 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_80_199 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_5855_ _5855_/A1 _6539_/A1 _5855_/B hold22/Z hold23/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi211_1
X_4806_ _7490_/Q _4809_/S _4807_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_119_121 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_119_110 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5786_ hold36/I _5520_/C _5786_/B1 _5792_/B1 _5786_/C1 _5802_/A1 _5787_/A3 VDD VSS
+ gf180mcu_fd_sc_mcu7t5v0__aoi222_1
X_4737_ hold467/Z _4748_/I1 _4741_/S _7453_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_147_452 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7525_ _7525_/D _7938_/RN _7961_/CLK _7525_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_175_783 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_174_282 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_174_260 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_7456_ _7456_/D _7877_/RN _7456_/CLK _7456_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
X_4668_ hold464/Z _3879_/Z _4668_/B hold465/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_134_124 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6407_ _4460_/Z _6417_/A2 _6407_/B _7832_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
Xhold930 hold930/I _4872_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
Xhold952 _7975_/Q _3632_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
Xhold963 _3768_/Z _7970_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
XFILLER_162_477 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_134_179 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_89_712 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7387_ _7387_/D _7938_/RN _7532_/CLK _7387_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
X_4599_ _4599_/A1 _6537_/A2 _4603_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
Xhold941 hold941/I _7551_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
X_6338_ hold682/Z _6349_/A2 _6339_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_104 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_89_778 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6269_ _4454_/Z _6281_/A2 _6269_/B _7767_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_48_108 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_8008_ _8008_/I _8008_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_84_494 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_71_100 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_56_196 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_71_144 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_44_32 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_13_712 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_40_531 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_40_553 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_157_227 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_100_71 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_12_277 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_138_463 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_60_64 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_166_794 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_125_124 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_4_443 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_140_105 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_153_499 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_140_116 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_79_211 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_69_73 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_95_759 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_67_428 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_94_247 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_47_141 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_47_152 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3970_ input49/Z _4275_/A2 _5886_/A1 input57/Z _4239_/A2 input25/Z _3998_/A2 VDD
+ VSS gf180mcu_fd_sc_mcu7t5v0__aoi222_1
X_5640_ _5640_/A1 _5520_/C _5640_/B1 _5640_/B2 _7541_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_31_564 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5571_ _5585_/A1 _5658_/B _5585_/B _5585_/C _5784_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XFILLER_79_2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_157_783 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_129_496 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4522_ _4522_/A1 _6537_/A2 _4526_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_7310_ _7900_/RN _4334_/Z _7310_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__and2_1
X_7241_ _7241_/A1 _7241_/A2 _7242_/C VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_4453_ hold11/Z _3810_/S hold12/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
Xhold226 hold226/I _7665_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
Xhold215 hold215/I _7739_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
Xhold204 _7611_/Q hold204/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
Xhold259 _7382_/Q hold259/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
Xhold237 _7819_/Q hold237/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
XFILLER_116_179 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xhold248 hold248/I _4496_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
X_4384_ _7511_/Q _7214_/A2 _7215_/C VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_98_531 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7172_ _7172_/A1 _7172_/A2 _7172_/A3 _7178_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand3_1
X_6123_ _6553_/A1 _6123_/A2 _6123_/B hold201/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
XTAP_531 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_520 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_542 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_140_672 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6054_ hold108/Z _6055_/A2 _6055_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_553 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_564 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_575 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_5005_ _3722_/I _3723_/I _5005_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__or2_2
XTAP_586 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_597 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_39_686 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_81_420 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1719 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_121_37 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1708 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_6956_ _7676_/Q _7191_/A2 _7204_/B1 _7766_/Q _6959_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_26_358 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_53_144 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5907_ _4454_/Z _5919_/A2 _5907_/B _7597_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_81_19 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_22_531 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6887_ _7469_/Q _6647_/Z _6887_/B1 _7510_/Q _6887_/C _6888_/A4 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi221_1
XFILLER_139_238 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_139_227 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5838_ _6547_/A1 _5840_/A2 _5838_/B _7567_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_22_586 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_155_709 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5769_ _5769_/A1 _5769_/A2 _5651_/Z _5769_/A4 _5770_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__and4_1
XFILLER_154_208 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_7508_ _7508_/D _7938_/RN _7532_/CLK _7508_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_107_124 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_107_113 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_30_34 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_146_34 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7439_ _7439_/D _7923_/RN _7599_/CLK _7988_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_30_67 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_135_499 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_116_680 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_89_531 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
Xhold771 _7393_/Q hold771/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
Xhold782 _7474_/Q hold782/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
Xhold760 hold760/I _7677_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
XFILLER_150_458 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
Xhold793 hold793/I _7534_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
XFILLER_39_10 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_49_406 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_162_33 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_89_597 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_49_428 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_130_193 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_76_247 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_29_141 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_44_122 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_32_328 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_13_553 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_158_536 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_158_525 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_40_383 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_139_783 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xoutput309 _8009_/Z spimemio_flash_io3_di VDD VSS gf180mcu_fd_sc_mcu7t5v0__buf_4
XFILLER_141_425 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_141_469 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_110_812 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_68_726 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_95_567 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_82_206 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_90_250 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6810_ _7804_/Q _6883_/A2 _6883_/B1 _7788_/Q _6812_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_63_464 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_35_144 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7790_ _7790_/D _7875_/RN _7790_/CLK _7790_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffsnq_1
XFILLER_177_812 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_149_514 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6741_ _7378_/Q _6882_/A2 _6880_/A2 _7817_/Q _6742_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_3953_ _3953_/A1 _3953_/A2 _3953_/A3 _3953_/A4 _3954_/A4 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand4_2
XFILLER_16_380 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_3884_ hold89/Z hold82/Z _6418_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_4
X_6672_ _7790_/Q _6893_/A2 _6659_/Z _7620_/Q _6673_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_176_333 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_137_709 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5623_ _5623_/A1 _5620_/B _5790_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_5554_ _5641_/A1 _5641_/A2 _5652_/A4 _5769_/A2 _5557_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand4_1
XFILLER_160_701 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_144_252 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5485_ _5680_/A1 _5779_/B1 _5485_/B _5504_/B1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_4505_ _4505_/A1 _6537_/A2 _4521_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_4
XFILLER_117_499 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_104_127 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_104_116 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7224_ _7224_/I0 _7945_/Q _7228_/S _7945_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_4436_ _7979_/Q _7875_/RN _4436_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__or2_1
X_4367_ _4367_/A1 _4367_/A2 _4367_/A3 _4372_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor3_1
XFILLER_160_756 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_132_458 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_116_37 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_104_149 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7155_ _7901_/Q _7197_/A2 _7195_/B1 _7627_/Q _7158_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_59_704 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6106_ _6553_/A1 _6106_/A2 _6106_/B hold189/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_101_812 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4298_ hold950/Z _4309_/S _4301_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_7086_ _7681_/Q _7191_/A2 _7190_/B1 _7617_/Q _7190_/A2 _7795_/Q _7089_/A2 VDD VSS
+ gf180mcu_fd_sc_mcu7t5v0__aoi222_1
XFILLER_86_545 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_86_534 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_372 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_394 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_383 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_6037_ hold190/Z _6038_/A2 _6038_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_39_450 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_39_461 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2217 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2206 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_92_18 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2239 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2228 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1505 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_12 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
X_7988_ _7988_/I _7988_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_1538 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1527 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1516 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_14_328 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_23 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_34 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_45 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_25_23 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_27_689 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_56 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_168_812 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1549 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_6939_ _6953_/A2 _6950_/A2 _6941_/A2 _7193_/C1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor3_4
XPHY_67 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_78 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_89 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_10_534 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_182_314 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_41_33 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_108_433 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_157_77 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_151_712 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xclkbuf_0_csclk _4416_/ZN clkbuf_0_csclk/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_123_425 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_9_2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xhold590 _7896_/Q hold590/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
XFILLER_2_744 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_150_266 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_110_108 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_89_361 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_77_523 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_49_203 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_173_98 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_77_567 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_66_63 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_66_52 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_18_601 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_49_269 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_17_144 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_18_656 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_72_272 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_72_250 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_159_812 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_32_136 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_173_314 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_158_388 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_127_753 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_154_550 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_5270_ _5292_/B _5624_/B _5391_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_5_582 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_114_458 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_99_169 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_99_158 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_87_309 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4221_ _7355_/Q _4488_/A1 _4554_/A1 _7385_/Q _4264_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_110_620 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_68_534 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4152_ hold609/Z _3963_/Z _4549_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_4083_ _7718_/Q hold90/I _4083_/B _4084_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_49_770 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7911_ _7911_/D _7923_/RN _7935_/CLK _7911_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffsnq_4
XFILLER_55_239 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_64_740 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_91_570 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7842_ _7842_/D _7901_/RN _7854_/CLK _7842_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_36_486 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_168_108 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4985_ _5022_/B _4943_/Z _5647_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_4
X_7773_ _7773_/D _7877_/RN _7773_/CLK _7773_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_63_283 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_24_659 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6724_ _7662_/Q _6885_/A2 _6644_/Z _7750_/Q _7776_/Q _6891_/C1 _6728_/A1 VDD VSS
+ gf180mcu_fd_sc_mcu7t5v0__aoi222_1
X_3936_ _3936_/A1 _3936_/A2 _3936_/A3 _3936_/A4 _3936_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__and4_1
X_3867_ _3886_/A2 hold54/Z _6248_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_4
X_6655_ _7910_/Q _6658_/A2 _6664_/A2 _6891_/B1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor3_4
X_3798_ hold49/Z hold52/Z _3800_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_5606_ _5735_/A2 _5658_/B _5752_/B1 _5606_/B _5610_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai31_1
XFILLER_118_742 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_118_720 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6586_ _6586_/A1 _6664_/A2 _6586_/B _6587_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_5537_ _5511_/C _5537_/A2 _5739_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_133_712 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_105_425 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_160_531 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_127_69 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5468_ _5031_/B _5473_/A2 _5471_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_7207_ _7961_/Q _7207_/A2 _7207_/B1 _7530_/Q _7207_/C _7208_/A4 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi221_1
XFILLER_160_575 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_5399_ _5735_/A2 _5585_/A1 _5724_/B _5759_/A1 _5735_/C _5401_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi221_1
X_4419_ _7979_/Q input88/Z _4420_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__or2_1
X_7138_ _7707_/Q _7190_/C1 _7196_/B1 _7643_/Q _7140_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_59_534 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_59_523 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7069_ _7778_/Q _7200_/A2 _7200_/B1 _7866_/Q _7075_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_59_567 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_100_174 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2025 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2014 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2003 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_100_196 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2058 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2047 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2036 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1313 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1302 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_54_250 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_55_773 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2069 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1357 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1346 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1335 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1324 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_15_637 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_42_423 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_146_2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1379 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1368 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_30_607 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_52_32 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_11_810 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_168_43 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_167_141 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xinput19 mask_rev_in[23] input19/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XFILLER_10_386 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_109_753 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_182_177 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_111_428 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_77_73 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_92_356 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_92_389 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_73_570 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_33_412 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_60_220 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_33_423 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1891 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1880 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_4770_ hold734/Z _4773_/A2 _4771_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_14_670 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_158_141 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3721_ _7908_/Q _6585_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__inv_1
XFILLER_174_656 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6440_ hold684/Z _6451_/A2 _6441_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_3652_ _7433_/Q _7001_/C VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_2
XFILLER_173_144 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_115_701 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_61_2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_6371_ _4454_/Z _6383_/A2 _6371_/B _7815_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_115_712 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_114_211 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5322_ _5689_/A2 _5687_/B _5724_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_2
XFILLER_142_531 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_142_575 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_114_266 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5253_ _5689_/A1 _5687_/B _5759_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_4
X_5184_ _5648_/A1 _5752_/B1 _5740_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_4204_ _4204_/A1 _4204_/A2 _4204_/A3 _4204_/A4 _7221_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor4_4
XFILLER_96_673 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4135_ hold42/Z hold149/Z _5841_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_3_70 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_29_718 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_113_16 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_83_312 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_83_301 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
Xclkbuf_leaf_63_csclk clkbuf_opt_1_0_csclk/Z _7738_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_56_526 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4066_ _7881_/Q _6503_/A1 _4488_/A1 _7358_/Q _6537_/A1 _7897_/Q _4067_/A4 VDD VSS
+ gf180mcu_fd_sc_mcu7t5v0__aoi222_1
XFILLER_24_401 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_36_250 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7825_ _7825_/D _7901_/RN _7873_/CLK _7825_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_24_445 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_36_272 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_169_428 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_24_467 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
Xclkbuf_leaf_78_csclk _7528_/CLK _7532_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_52_765 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4968_ _5006_/B _5254_/A2 _5709_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_4
X_7756_ _7756_/D _7875_/RN _7830_/CLK _7756_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_51_286 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_4899_ _5006_/B _5006_/C _5392_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_2
XFILLER_149_163 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_149_141 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7687_ _7687_/D _7923_/RN _7698_/CLK _7687_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
X_3919_ _4284_/A1 _7230_/A1 _3921_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_6707_ _6707_/A1 _6767_/C _6707_/B1 _6707_/B2 _7433_/Q _6708_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi221_1
XFILLER_20_662 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_20_673 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6638_ _6878_/A2 _6658_/A2 _6664_/A2 _6893_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor3_4
XFILLER_165_667 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_138_57 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_138_46 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_106_734 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6569_ _7435_/Q _6622_/A2 _6569_/A3 _6571_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor3_1
XFILLER_133_553 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xclkbuf_leaf_16_csclk _7873_/CLK _7869_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_154_34 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_120_203 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_154_56 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_120_247 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_93_109 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_86_172 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_170_66 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_74_334 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_47_87 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_74_389 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_34_209 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_55_570 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_103_93 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1121 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1132 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1110 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_15_423 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_27_283 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1165 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1154 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1143 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1198 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1187 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1176 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_43_798 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_156_601 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_8_37 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_7_633 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_7_622 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_7_611 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_156_689 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_156_656 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_155_144 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_143_306 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_128_347 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_109_550 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_7_655 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_171_637 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_109_561 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_6_176 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_124_531 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_905 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_916 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_88_83 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_927 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_938 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_949 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_111_247 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_78_673 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_78_695 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_92_164 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_92_153 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_18_250 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_5940_ hold885/Z _5953_/A2 _5941_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_92_197 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_179_737 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7610_ _7610_/D _7923_/RN _7820_/CLK _7610_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_21_404 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5871_ _5871_/A1 _6537_/A2 _5873_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_178_247 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_33_286 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4822_ _7498_/Q _4828_/S _4823_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_4753_ hold263/Z _4753_/I1 _4753_/S _4753_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_7541_ _7541_/D _7959_/RN _7545_/CLK hold40/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
X_3704_ _7671_/Q _3704_/ZN VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_7472_ _7472_/D _7961_/RN _7531_/CLK _7472_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
X_4684_ _7465_/Q _3879_/Z _4684_/B _4685_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_107_509 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6423_ hold671/Z _6434_/A2 _6424_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_3635_ _3635_/I _3958_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_6354_ _4454_/Z _6366_/A2 _6354_/B _7807_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_108_27 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_170_670 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5305_ _5682_/A1 _5692_/A2 _5307_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_6285_ hold877/Z _6298_/A2 _6286_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_5236_ _5200_/B _3727_/I _5421_/A1 _5621_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__and3_2
XFILLER_130_534 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_115_597 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_88_459 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_124_37 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_102_258 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_102_247 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_69_651 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_5167_ _5735_/A2 _5672_/A2 _5167_/B _5171_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_124_48 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_56_323 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5098_ _5098_/A1 _5098_/A2 _5772_/A1 _5749_/A1 _5106_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand4_1
X_4118_ _4141_/A1 _3963_/Z _4853_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_4049_ _4049_/A1 _4049_/A2 _4058_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_84_676 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_17_35 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_37_570 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_56_389 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_215 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_204 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_169_225 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7808_ _7808_/D _7877_/RN _7812_/CLK _7808_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffsnq_1
XPHY_259 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_248 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_237 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_226 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_25_798 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_178_770 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7739_ _7739_/D _7923_/RN _7816_/CLK _7739_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_137_122 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_137_144 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_165_486 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_153_626 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_153_637 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_137_177 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_125_306 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_165_33 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_152_147 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_109_2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_106_531 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_121_578 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_121_567 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_58_64 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xhold8 hold8/I hold8/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
XFILLER_114_92 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_90_602 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_74_63 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_16_721 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_15_242 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_15_286 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_70_392 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_143_103 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
Xhold408 _7509_/Q hold408/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
Xhold419 _4749_/Z _7462_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
XFILLER_7_496 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_98_724 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_112_534 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_97_212 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_713 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_702 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_724 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_6070_ _4481_/I _6072_/A2 _6070_/B hold512/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
XTAP_735 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_746 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_757 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_768 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_5021_ _5529_/A2 _5529_/A3 _5021_/B1 _5010_/Z _5548_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_4
XFILLER_24_2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_779 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_66_632 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_66_676 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_65_153 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_26_529 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_38_356 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_38_389 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_80_134 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6972_ _7798_/Q _7191_/B1 _7201_/B1 _7668_/Q _6972_/C _6976_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi221_1
XFILLER_19_570 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_53_337 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_110_17 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5923_ hold883/Z _5936_/A2 _5924_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_5854_ _7982_/I _5855_/A1 _5855_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_21_212 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_179_567 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_166_206 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_21_223 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4805_ _7224_/I0 _7489_/Q _4809_/S _7489_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_119_100 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5785_ _5785_/A1 _5795_/A3 _5785_/A3 _5785_/B _5787_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai31_1
X_7524_ _7524_/D _7938_/RN _7639_/CLK _7524_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
X_4736_ hold34/Z hold32/Z _4741_/S hold35/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_119_144 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_174_272 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_174_250 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4667_ _3879_/Z hold64/I _4668_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_7455_ _7455_/D _7853_/RN _7600_/CLK _7455_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_135_615 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_119_155 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6406_ hold683/Z _6417_/A2 _6407_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
Xhold920 hold920/I _6094_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
Xhold931 hold931/I _7528_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
X_7386_ _7386_/D _7875_/RN _7822_/CLK _7386_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
Xhold964 hold11/I hold964/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
Xhold953 _7339_/Q hold953/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
XFILLER_115_361 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6337_ _4454_/Z _6349_/A2 _6337_/B _7799_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_4598_ _4454_/Z _4598_/A2 _4598_/B _7402_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
Xhold942 _7548_/Q hold942/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
XFILLER_143_692 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_135_25 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_103_567 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6268_ hold901/Z _6281_/A2 _6269_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_5219_ _5452_/C _5543_/C _5545_/A2 _5580_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor3_2
XFILLER_130_364 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6199_ hold128/Z _6208_/A2 hold129/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_8007_ _8007_/I _8007_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_28_23 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_28_34 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_72_602 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_57_687 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_52_392 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_138_420 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_8_205 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_166_751 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_165_283 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_5_16 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_4_433 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_180_264 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_109_81 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_109_70 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_79_223 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_48_632 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_85_73 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_63_602 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_48_676 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_51_808 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_50_318 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_176_504 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5570_ _5692_/A1 _5218_/C _5702_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_156_250 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_144_401 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_116_103 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4521_ _6553_/A1 _4521_/A2 _4521_/B hold359/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_4452_ hold49/Z hold567/Z _4455_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_7240_ _7520_/Q _7240_/A2 _7240_/B1 _7519_/Q _7241_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_1
Xhold216 _7970_/Q hold216/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
XFILLER_171_220 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
Xhold205 hold205/I _5936_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
Xhold227 _7729_/Q hold227/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
Xhold238 hold238/I _7819_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
Xhold249 hold249/I _7358_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
XFILLER_171_286 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4383_ _4383_/A1 _4383_/A2 _4383_/B _7413_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_7171_ _7527_/Q _7189_/A2 _7191_/B1 _7405_/Q _7172_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_6122_ hold199/Z _6123_/A2 hold200/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_543 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_532 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_521 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_510 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_6053_ hold233/Z _6055_/A2 _6053_/B _7666_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_105_39 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_105_17 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_86_727 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_85_215 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_554 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_565 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_576 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_5004_ _3722_/I _3723_/I _5254_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_4
XTAP_587 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_598 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_38_120 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_54_602 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_93_292 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_26_315 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_39_698 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1709 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_6955_ _7914_/Q _7913_/Q _6599_/Z _6955_/A4 _7205_/B1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor4_4
XFILLER_53_156 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5906_ hold615/Z _5919_/A2 _5907_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_179_364 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_34_392 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6886_ _6886_/A1 _6886_/A2 _6886_/A3 _6887_/C VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_179_386 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_10_727 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5837_ hold647/Z _5840_/A2 _5838_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_22_576 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5768_ _5122_/Z _5768_/A2 _5768_/A3 _5769_/A4 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_175_570 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4719_ _4719_/A1 _6537_/A2 _4731_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_4
X_7507_ _7507_/D _7938_/RN _7532_/CLK _7507_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_147_283 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5699_ _5590_/B _5581_/B _5737_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_7438_ _7438_/D _7923_/RN _7597_/CLK _7438_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_107_169 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_107_158 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_163_798 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
Xhold761 _7996_/I hold761/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
X_7369_ _7369_/D _7875_/RN _7567_/CLK _7369_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffsnq_1
XFILLER_1_425 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xhold772 _7558_/Q hold772/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
Xhold750 _7387_/Q hold750/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
Xhold794 _7790_/Q hold794/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
Xhold783 _7782_/Q hold783/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
XFILLER_45_602 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_57_462 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_176_2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_44_112 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_57_473 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_60_605 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_32_318 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_138_250 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_138_283 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_138_272 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_126_445 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_181_540 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_126_456 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_181_595 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_153_286 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_113_128 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_113_117 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_99_329 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_122_673 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_67_215 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_96_72 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_95_546 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_36_602 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_48_495 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6740_ _7719_/Q _6881_/A2 _6882_/B1 _7655_/Q _6742_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_50_104 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_51_638 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3952_ _7738_/Q _6192_/A1 _6090_/A1 _7690_/Q _3953_/A4 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_16_392 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_3883_ _3886_/A2 _4075_/B _4232_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_4
XFILLER_91_2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6671_ _7814_/Q _6880_/A2 _6892_/A2 _7758_/Q _6673_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_5622_ _5622_/A1 _5620_/B _5622_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__or2_1
XFILLER_176_389 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_157_570 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_5553_ _5553_/A1 _5553_/A2 _5769_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_129_294 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_129_283 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4504_ _6553_/A1 _4504_/A2 _4504_/B hold362/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_5484_ _4965_/B _5603_/A1 _5797_/A2 _5485_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor3_1
XFILLER_145_798 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_132_415 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7223_ _7223_/A1 _7228_/S _7223_/B _7944_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_4435_ _7980_/Q _7875_/RN _4435_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__or2_1
X_4366_ _4366_/A1 _4366_/A2 _4367_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_7154_ _7651_/Q _7195_/A2 _7207_/B1 _7723_/Q _7158_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_6105_ hold187/Z _6106_/A2 hold188/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_100_301 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_4297_ _7342_/Q _4308_/S _4296_/Z _4297_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__and3_1
XFILLER_112_194 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7085_ _7705_/Q _7190_/C1 _7089_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_373 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_384 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_132_15 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_67_760 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6036_ _4481_/I _6038_/A2 _6036_/B _7658_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
XTAP_395 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2207 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_132_37 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_100_389 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2229 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2218 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1506 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_82_741 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_13 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
X_7987_ _7987_/I _7987_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_1539 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1528 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1517 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_14_318 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_24 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_35 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_46 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_25_13 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_25_35 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_42_605 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_54_498 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_155_7 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6938_ _6938_/I _6948_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XPHY_57 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_68 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_79 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_179_172 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6869_ _7509_/Q _6887_/B1 _6891_/B1 _7507_/Q _6871_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_182_326 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_150_212 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_135_286 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_123_437 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_151_768 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
Xhold580 hold580/I hold580/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
XFILLER_150_278 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_104_673 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xhold591 hold591/I _6543_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
XFILLER_49_215 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_18_646 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_45_443 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_32_104 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_33_638 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_60_479 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_158_334 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_13_384 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_173_304 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_139_570 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_9_366 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_40_192 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_63_6 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_141_212 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_5_561 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_141_245 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_99_148 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4220_ _7766_/Q _6265_/A1 _4564_/A1 _7389_/Q _4264_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_4151_ hold609/Z _4151_/A2 _4888_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_110_676 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_95_354 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4082_ _7726_/Q hold28/I _6124_/A1 _7702_/Q _4084_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_7910_ _7910_/D _7938_/RN _7940_/CLK _7910_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffsnq_4
X_7841_ _7841_/D _7901_/RN _7899_/CLK _7841_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_64_730 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_63_273 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_24_605 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4984_ _3723_/I _5777_/A1 _5797_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_2
X_7772_ _7772_/D _7901_/RN _7866_/CLK _7772_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
X_6723_ _7784_/Q _6883_/B1 _6894_/A2 _7840_/Q _6729_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_3935_ input27/Z _4239_/A2 _6537_/A1 _7900_/Q _3936_/A4 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_51_479 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_20_811 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6654_ _6878_/A2 _6658_/A2 _6662_/A3 _6891_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor3_4
XFILLER_137_507 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_109_209 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5605_ _5735_/A2 _5606_/B _5674_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_3866_ hold54/Z _3847_/Z _6265_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_4
X_3797_ _7341_/Q _7414_/Q _4303_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_6585_ _7909_/Q _6585_/A2 _6664_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_4
X_5536_ _5543_/B _5153_/C _5536_/A3 _5537_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor3_1
XFILLER_145_562 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_118_765 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_133_724 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_132_212 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5467_ _5602_/A1 _5602_/A2 _5527_/A1 _5473_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor3_1
XFILLER_117_286 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_105_415 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_172_392 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_127_59 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_105_459 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4418_ input83/Z _4418_/I1 _7979_/Q _4418_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_7206_ _7206_/A1 _7206_/A2 _7206_/A3 _7207_/C VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_99_682 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5398_ _5733_/A2 _5398_/A2 _5586_/A3 _5398_/A4 _5414_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand4_1
X_7137_ _7675_/Q _7201_/B1 _7204_/B1 _7773_/Q _7140_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_98_181 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_86_321 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_59_546 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_4349_ _7902_/Q _6565_/A1 _6622_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_143_69 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7068_ _7068_/A1 _7068_/A2 _7068_/A3 _7068_/A4 _7078_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand4_1
XFILLER_86_387 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_74_538 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6019_ _4481_/I _6021_/A2 _6019_/B _7650_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
XTAP_2015 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2004 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_36_34 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_55_730 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2059 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2048 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2026 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2037 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1314 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1303 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1347 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1336 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1325 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_70_744 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_15_649 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1358 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1369 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_23_682 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_168_676 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_139_2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_10_321 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_170_318 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_123_212 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_2_531 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_151_587 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_117_70 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_78_811 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_2_575 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_77_354 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_77_96 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_77_85 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_93_73 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_93_62 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1870 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_60_254 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_33_468 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1892 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1881 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_61_799 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_3720_ _7909_/Q _6636_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__inv_1
XFILLER_174_602 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_9_141 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_174_646 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_146_326 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_3651_ _7905_/Q _6571_/B2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_146_348 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6370_ hold915/Z _6383_/A2 _6371_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_5321_ _5724_/B _5648_/B2 _5496_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_114_201 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_54_2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_154_392 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_142_521 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5252_ _5199_/B _5201_/B _3728_/I _5022_/B _5687_/C VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand4_4
X_5183_ _5496_/A1 _5099_/B _5512_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_68_321 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4203_ _4203_/A1 _4203_/A2 _4203_/A3 _4203_/A4 _4204_/A4 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand4_2
X_4134_ hold149/Z _3869_/I _4754_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_56_505 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_83_357 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4065_ _7817_/Q _6367_/A1 hold150/I _7566_/Q _4231_/B1 input67/Z _4067_/A3 VDD VSS
+ gf180mcu_fd_sc_mcu7t5v0__aoi222_1
X_7824_ _7824_/D _7901_/RN _7896_/CLK _7824_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffsnq_1
XFILLER_91_390 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_51_221 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_52_744 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7755_ hold7/Z _7877_/RN _7755_/CLK _7755_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
X_4967_ _3722_/I _3723_/I _5206_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_4
X_4898_ _5006_/B _5006_/C _4898_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__and2_2
X_3918_ _3918_/A1 _3918_/A2 _3917_/Z _7230_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor3_4
X_7686_ _7686_/D _7923_/RN _7734_/CLK _7686_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffsnq_1
X_6706_ _6706_/A1 _6706_/A2 _6706_/A3 _6707_/B2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor3_1
X_3849_ hold42/Z _4141_/A1 _6073_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_4
X_6637_ _7910_/Q _6661_/A3 _6658_/A3 _6880_/C2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor3_4
XFILLER_180_605 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_22_69 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6568_ _7904_/Q _6561_/Z _6570_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_5519_ _5519_/A1 _5519_/A2 _5519_/B _5520_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_152_318 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_98_18 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_105_212 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xclkbuf_3_2__f_csclk clkbuf_0_csclk/Z _7528_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
X_6499_ hold664/Z _6502_/A2 _6500_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_133_565 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_79_608 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_87_641 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_59_354 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_47_505 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_170_45 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_170_34 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_47_99 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_70_530 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1122 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1111 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1100 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_28_796 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_43_733 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_43_722 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_179_10 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1155 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1144 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1133 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1199 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1188 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1177 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1166 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_15_479 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_30_427 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_30_438 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_42_276 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_168_451 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_11_641 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_30_449 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_128_315 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_109_584 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_170_137 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_136_392 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_88_62 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_906 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_917 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_151_373 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_111_215 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_97_438 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_97_449 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_928 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_939 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_120_760 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_93_600 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_65_357 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_92_176 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_92_143 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_19_763 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_53_519 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5870_ _5870_/A1 hold47/Z _5870_/B hold22/Z hold48/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XFILLER_34_744 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4821_ _7221_/A1 _4828_/S _4821_/B _7497_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_34_755 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2390 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_61_596 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_61_585 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_61_574 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4752_ _4481_/I _4753_/S _4752_/B _7464_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_7540_ _7540_/D _7959_/RN _7545_/CLK hold74/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_21_438 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4683_ _3879_/Z hold2/Z _4684_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_3703_ _7679_/Q _3703_/ZN VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_7471_ _7471_/D _7961_/RN _7627_/CLK _7471_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_162_605 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_146_123 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_135_808 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3634_ _3634_/I _4402_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_6422_ _4454_/Z _6434_/A2 _6422_/B _7839_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_162_627 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_134_318 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_108_17 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6353_ hold830/Z _6366_/A2 _6354_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_5304_ _5319_/B _5692_/A2 _5307_/B2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_103_716 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6284_ _6539_/A1 _6298_/A2 _6284_/B _7774_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_5235_ _5685_/B _5292_/B _5614_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_69_641 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5166_ _5643_/A2 _5783_/A2 _5166_/B _5166_/C _5171_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XFILLER_96_460 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_84_622 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_56_313 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5097_ _5735_/A2 _5669_/A1 _5749_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_4117_ hold54/Z _3959_/Z _4574_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_71_305 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4048_ input55/Z _5886_/A1 _4239_/A2 input23/Z _5870_/A1 _7576_/Q _4049_/A2 VDD VSS
+ gf180mcu_fd_sc_mcu7t5v0__aoi222_1
XFILLER_140_37 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_169_215 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_216 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_205 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_40_703 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_7807_ _7807_/D _7877_/RN _7809_/CLK _7807_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffsnq_1
XPHY_249 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_238 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_227 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
X_5999_ hold724/Z _6004_/A2 _6000_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_24_276 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7738_ _7738_/D _7938_/RN _7738_/CLK _7738_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_33_35 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_40_747 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_149_57 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_20_460 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_138_646 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_20_471 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7669_ _7669_/D _7938_/RN _7791_/CLK _7669_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffsnq_1
XFILLER_165_476 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_153_649 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_118_392 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_106_598 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_106_587 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
Xoutput290 _7366_/Q pll_trim[3] VDD VSS gf180mcu_fd_sc_mcu7t5v0__buf_4
Xhold9 hold9/I hold9/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
XFILLER_75_600 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_59_140 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_101_281 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_74_132 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_59_195 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_63_806 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_47_357 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_74_187 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_74_176 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_74_53 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_62_338 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_15_232 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_15_221 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_31_736 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_43_574 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_90_41 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_30_246 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_90_74 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_144_605 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_116_318 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xclkbuf_leaf_62_csclk clkbuf_3_6__f_csclk/Z _7736_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
Xhold409 _7494_/Q hold409/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
XFILLER_171_479 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_152_671 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_98_747 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xclkbuf_leaf_77_csclk _7528_/CLK _7531_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XTAP_714 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_703 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_725 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_5020_ _5010_/Z _5021_/B1 _5020_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_97_235 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_736 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_747 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_758 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_78_471 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_78_460 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_769 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_17_2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_38_379 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_93_496 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_81_625 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_81_636 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_80_124 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6971_ _6971_/A1 _6971_/A2 _6971_/A3 _6972_/C VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_0_50 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_72 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5922_ hold47/Z _5936_/A2 _5922_/B hold502/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_5853_ hold50/Z hold106/Z _5853_/S _5853_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
Xclkbuf_leaf_15_csclk _7873_/CLK _7901_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_80_179 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5784_ _5784_/A1 _5704_/Z _5784_/A3 _5785_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_22_747 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4804_ _7223_/A1 _4809_/S _4804_/B _7488_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_175_730 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4735_ _7451_/Q hold13/Z _4741_/S hold14/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_147_421 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_9_70 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7523_ _7523_/D _7938_/RN _7606_/CLK _7523_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
X_4666_ _7984_/I _4685_/A1 _4669_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_7454_ _7454_/D _7853_/RN _7600_/CLK _7454_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_119_178 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_119_38 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_135_638 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xhold921 hold921/I _7685_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
X_4597_ hold833/Z _4598_/A2 _4598_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_7385_ _7385_/D _7875_/RN _7547_/CLK _7385_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
Xhold910 _7669_/Q hold910/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
X_6405_ _4454_/Z _6417_/A2 _6405_/B _7831_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
Xhold943 _7954_/Q _3671_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
Xhold954 _7977_/Q _3745_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
X_6336_ hold875/Z _6349_/A2 _6337_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
Xhold932 _7553_/Q _3636_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
Xhold965 hold30/I hold965/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
XFILLER_143_682 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_115_384 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_1_629 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_130_321 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_95_19 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_139 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6267_ _6539_/A1 _6281_/A2 _6267_/B _7766_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_5218_ _5421_/B1 _5218_/A2 _5218_/B _5218_/C _5294_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai211_1
X_6198_ _4460_/Z _6208_/A2 _6198_/B hold640/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_8006_ _8006_/I _8006_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_29_302 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_57_600 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5149_ _5543_/B _5552_/A3 _5548_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_97_791 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_84_463 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_29_357 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_29_379 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_45_806 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_84_496 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_56_176 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_44_34 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_13_703 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_44_67 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_13_769 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_153_402 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_138_476 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_126_605 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_125_104 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_121_2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_176_99 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_125_126 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_5_28 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_153_479 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_125_148 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_106_384 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_4_489 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_69_97 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_684 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_90_422 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_90_411 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_75_496 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_47_198 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_62_179 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_62_168 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_149_708 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_31_544 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_129_421 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_79_4 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_157_774 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_11_290 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4520_ hold357/Z _4521_/A2 hold358/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_172_733 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
Xhold217 hold217/I _4476_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
XFILLER_156_273 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_117_638 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xhold206 hold206/I _7611_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
X_4451_ hold927/Z _4487_/A1 _4456_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_7_283 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xhold228 hold228/I _7729_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
XFILLER_144_457 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xhold239 _7869_/Q hold239/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
X_7170_ _7521_/Q _7189_/B1 _7189_/C1 _7494_/Q _7172_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_4382_ _4383_/A2 _4382_/A2 _7413_/Q _4383_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_6121_ _4481_/I _6123_/A2 _6121_/B hold703/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
XTAP_500 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_112_321 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_98_566 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_98_555 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_98_544 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_533 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_522 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_511 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_6052_ hold392/Z _6055_/A2 _6053_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_86_717 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_544 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_555 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_566 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_5003_ _5087_/C _5777_/A1 _5741_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_2
XTAP_577 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_588 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_599 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_66_463 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_38_176 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6954_ _6955_/A4 _6954_/A2 _7205_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_4
X_5905_ hold47/Z _5919_/A2 _5905_/B hold369/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_81_499 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_179_354 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6885_ _7505_/Q _6885_/A2 _6885_/B1 _7528_/Q _6886_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_14_37 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_5836_ _6545_/A1 _5840_/A2 _5836_/B hold151/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_5767_ _5331_/Z _5767_/A2 _5767_/A3 _5771_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand3_1
X_7506_ _7506_/D _7959_/RN _7959_/CLK hold49/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_4
X_4718_ _4718_/A1 _4718_/A2 _4718_/B hold133/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_5698_ _5684_/Z _5698_/A2 _5698_/B _5719_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_108_605 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4649_ hold323/Z _4652_/A1 hold324/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_107_115 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7437_ _7437_/D _7923_/RN _7597_/CLK _7437_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_163_766 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
Xhold762 hold762/I _7422_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
XFILLER_150_416 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
Xhold740 _7998_/I hold740/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
Xhold773 _7563_/Q hold773/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
XFILLER_1_415 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_7368_ _7368_/D _7961_/RN _7570_/CLK _7368_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffsnq_1
Xhold751 _7582_/Q hold751/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
X_7299_ _7901_/RN _4334_/Z _7299_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_131_641 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xhold784 _7798_/Q hold784/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
Xhold795 _7846_/Q hold795/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
XFILLER_1_437 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6319_ hold925/Z _6332_/A2 _6320_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_103_354 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_85_783 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_55_33 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_169_2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_45_658 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_72_477 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_44_179 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_111_83 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_71_98 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_166_593 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_154_744 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_153_232 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_5_754 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_122_630 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_95_503 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_95_558 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_83_709 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_492 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_48_463 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_91_753 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_35_146 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3951_ _7714_/Q _6141_/A1 hold90/I _7722_/Q _3953_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_63_499 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_50_138 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3882_ _4075_/B _3881_/Z _4219_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_4
X_6670_ _7644_/Q _6880_/C2 _6644_/Z _7748_/Q _6673_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_5621_ _5624_/A2 _5648_/B2 _5621_/B _5740_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_84_2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5552_ _5543_/B _5153_/C _5552_/A3 _5552_/A4 _5553_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor4_1
XFILLER_157_582 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_129_273 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_4503_ hold360/Z _4504_/A2 hold361/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_5483_ _5543_/C _5543_/B _5498_/A2 _5498_/B _5218_/B _5547_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai32_1
X_4434_ _7520_/Q _4338_/Z _7512_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__and2_1
X_7222_ _7944_/Q _7228_/S _7223_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_4365_ _5224_/A3 _5224_/A4 _4365_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__or2_1
XFILLER_160_747 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_113_641 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7153_ _7153_/A1 _7153_/A2 _7153_/A3 _7153_/A4 _7159_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand4_1
XFILLER_140_460 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_101_803 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7084_ _7753_/Q _7201_/A2 _7201_/B1 _7673_/Q _7100_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_6104_ _4481_/I _6106_/A2 _6104_/B hold707/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_4296_ _7341_/Q _7340_/Q _4296_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_86_547 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6035_ hold509/Z _6038_/A2 _6036_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_374 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_385 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_58_238 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_396 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2208 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_82_720 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_73_219 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_67_783 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_67_772 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_39_496 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2219 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_82_731 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_15_809 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_26_124 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_162_9 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1529 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1518 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1507 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_7986_ _7986_/I _7986_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XPHY_25 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_14 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_36 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_47 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_26_179 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_41_105 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_42_617 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6937_ _6937_/A1 _6954_/A2 _6938_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_4
XPHY_58 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_69 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
X_6868_ _7470_/Q _6659_/Z _6884_/B1 _7521_/Q _6871_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_41_149 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_167_357 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_10_514 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5819_ _6539_/A1 _5827_/A2 _5819_/B _7558_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_6799_ _6799_/A1 _6799_/A2 _6799_/A3 _6799_/A4 _6799_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__and4_1
XFILLER_41_35 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_182_349 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_136_733 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_157_79 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xhold570 hold570/I _7417_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
XFILLER_173_34 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_1_212 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xhold581 hold581/I _7571_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
Xhold592 hold592/I _7896_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
XFILLER_2_18 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_65_709 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_72_263 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_26_691 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_45_499 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_13_352 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_158_346 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_9_378 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_154_530 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_181_371 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_127_799 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_126_276 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_114_405 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_142_758 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_142_747 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_122_460 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_110_600 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_96_812 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4150_ hold38/Z _4217_/A2 _4848_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_4081_ _7734_/Q _6192_/A1 _6073_/A1 _7678_/Q _6107_/A1 _7694_/Q _4084_/A1 VDD VSS
+ gf180mcu_fd_sc_mcu7t5v0__aoi222_1
XFILLER_64_720 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_49_783 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_102_19 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_7840_ _7840_/D _7901_/RN _7864_/CLK _7840_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffsnq_1
XFILLER_64_753 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_36_444 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4983_ _5206_/A2 _5709_/A1 _5669_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_4
X_7771_ _7771_/D _7877_/RN _7873_/CLK _7771_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_51_436 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_51_447 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_177_611 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6722_ _7377_/Q _6882_/A2 _6712_/Z _6830_/B _6894_/C1 _7832_/Q _6729_/A2 VDD VSS
+ gf180mcu_fd_sc_mcu7t5v0__aoi222_1
X_3934_ _7381_/Q hold55/I _4505_/A1 _7369_/Q _6452_/A1 _7860_/Q _3936_/A3 VDD VSS
+ gf180mcu_fd_sc_mcu7t5v0__aoi222_1
X_3865_ _4212_/A2 hold149/Z _5920_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_4
XFILLER_32_672 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_32_683 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6653_ _6878_/A2 _6663_/A4 _6662_/A3 _6890_/B1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor3_4
XFILLER_149_357 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_5604_ _4943_/Z _5604_/A2 _5606_/B _5610_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_176_176 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_164_327 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3796_ _3783_/Z _3925_/A2 hold75/I hold71/Z hold72/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__or4_4
X_6584_ _6587_/A2 _6584_/A2 _7908_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_5535_ _5535_/A1 _5548_/A3 _5536_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_118_755 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_118_744 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_11_27 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5466_ _5735_/A2 _4996_/Z _5658_/B _5643_/A2 _5674_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_4417_ input84/Z input67/Z _7980_/Q _4417_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_7205_ _7534_/Q _7205_/A2 _7205_/B1 _7538_/Q _7206_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_120_408 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_5397_ _5669_/B _5669_/A1 _5292_/B _5621_/B _5583_/B _5398_/A4 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi221_1
XFILLER_160_599 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_141_780 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_99_694 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7136_ _7781_/Q _7200_/A2 _7203_/B1 _7885_/Q _7140_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_98_171 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_98_160 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_59_536 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4348_ _7902_/Q _6565_/A1 _6622_/A1 _7581_/Q _6572_/A1 _7432_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai32_1
X_7067_ _7712_/Q _7189_/A2 _7189_/B1 _7688_/Q _7189_/C1 _7656_/Q _7068_/A4 VDD VSS
+ gf180mcu_fd_sc_mcu7t5v0__aoi222_1
XFILLER_47_709 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4279_ _4279_/A1 _4279_/A2 _4279_/A3 _4279_/A4 _4279_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__and4_1
XFILLER_100_176 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_74_528 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6018_ hold659/Z _6021_/A2 _6019_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_46_208 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2016 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2005 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_27_422 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_27_444 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_160_6 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2049 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2038 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2027 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1304 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_7969_ _7969_/D _7322_/Z _7972_/CLK hold15/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XTAP_1348 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1337 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1326 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1315 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_14_105 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_15_628 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_27_499 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_42_425 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1359 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_11_812 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_52_34 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_168_34 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_156_806 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_109_700 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_167_176 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_182_168 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_108_276 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_108_254 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_124_747 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_151_566 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_96_108 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_117_82 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_104_460 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_133_70 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_46_753 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_92_369 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_61_712 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_61_701 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_18_455 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_93_85 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_33_425 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_159_611 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1860 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_61_778 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1893 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1882 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1871 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_20_108 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_158_143 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_13_171 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_158_176 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3650_ _7904_/Q _6567_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_161_308 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5320_ _5006_/C _5419_/B _5555_/B _5326_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_5251_ _5338_/A1 _5369_/B _5271_/A3 _5624_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor3_4
XFILLER_102_419 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_69_812 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4202_ _4202_/A1 _4202_/A2 _4202_/A3 _4203_/A4 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor3_1
XFILLER_47_2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5182_ _5797_/B _5797_/C _5741_/A3 _5185_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor3_1
XFILLER_123_780 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_95_141 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_3_83 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_29_709 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4133_ _4141_/A1 _4155_/A2 _4858_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_2
XFILLER_110_463 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4064_ _7607_/Q _5920_/A1 _4505_/A1 _7366_/Q _6005_/A1 hold78/I _4067_/A2 VDD VSS
+ gf180mcu_fd_sc_mcu7t5v0__aoi222_1
XFILLER_95_185 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_37_731 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_64_550 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_7823_ _7823_/D _7875_/RN _7823_/CLK _7823_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffsnq_1
X_7754_ _7754_/D _7877_/RN _7755_/CLK _7754_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_24_458 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_24_469 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_149_121 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4966_ _5309_/A1 _5087_/C _4969_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_6705_ _6705_/A1 _6705_/A2 _6705_/A3 _6705_/A4 _6706_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand4_1
X_3917_ _3917_/A1 _3917_/A2 _3917_/A3 _3917_/A4 _3917_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__or4_1
X_7685_ _7685_/D _7923_/RN _7815_/CLK _7685_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffsnq_1
X_4897_ _4454_/Z _4897_/A2 _4897_/B hold798/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_177_496 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_165_636 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_149_176 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_149_165 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3848_ _4141_/A1 _3847_/Z _6141_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_4
XFILLER_22_37 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_6636_ _6636_/A1 _7908_/Q _6658_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_4
X_3779_ _7977_/Q hold936/Z _3780_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_138_37 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_4_808 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6567_ _6567_/A1 _6565_/B _6567_/B1 _6557_/I _7904_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai22_1
XFILLER_164_179 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5518_ _5547_/A1 _5518_/A2 _5518_/A3 _5519_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor3_1
XFILLER_106_747 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6498_ _6549_/A1 _6502_/A2 _6498_/B _7875_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_5449_ _5714_/A1 _5797_/A2 _5543_/C _5452_/C _5450_/C VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XFILLER_78_108 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_160_396 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_121_728 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_7119_ _7650_/Q _7195_/A2 _7195_/B1 _7626_/Q _7195_/C1 _7876_/Q _7121_/A3 VDD VSS
+ gf180mcu_fd_sc_mcu7t5v0__aoi222_1
XFILLER_59_366 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_47_34 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_47_517 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_47_528 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_101_496 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_103_73 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_1123 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1112 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1101 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_63_22 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_15_425 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_43_712 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_55_583 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
Xclkbuf_1_1__f_wbbd_sck clkbuf_0_wbbd_sck/Z net299_2/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_151_2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_103_95 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1156 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1145 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1134 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_244 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1189 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1178 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1167 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_70_597 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_42_266 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_168_463 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_168_441 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_129_806 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_8_17 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_7_624 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_11_697 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_10_185 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_6_134 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_170_105 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_155_157 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_164_680 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_109_596 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_112_717 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_907 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_105_791 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_105_780 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_97_428 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_88_85 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_918 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_929 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_77_141 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_92_155 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_81_807 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_19_775 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_34_734 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_2380 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_179_739 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4820_ _7497_/Q _4828_/S _4821_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_2391 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_21_428 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4751_ hold520/Z _4753_/S _4752_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_1
XTAP_1690 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_174_422 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_159_496 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_147_636 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4682_ hold229/Z _4685_/A1 hold230/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_3702_ _7687_/Q _3702_/ZN VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_7470_ _7470_/D _7961_/RN _7531_/CLK _7470_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
X_3633_ _7973_/Q _3765_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_6421_ hold872/Z _6434_/A2 _6422_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_146_179 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6352_ hold47/Z _6366_/A2 _6352_/B _7806_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_142_330 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5303_ _3728_/I _5022_/B _5303_/A3 _5303_/A4 _5692_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand4_4
XFILLER_103_706 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6283_ hold786/Z _6298_/A2 _6284_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_5234_ _5687_/B _5365_/B1 _5292_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_4
XFILLER_88_428 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5165_ _5006_/B _5206_/A2 _5476_/B _5319_/C _5692_/B _5645_/A1 _5166_/C VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai33_1
XFILLER_124_17 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_111_783 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_111_772 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_4116_ hold54/Z _3963_/Z _4522_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_5096_ _5669_/A1 _5783_/A2 _5772_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_4047_ _7378_/Q hold55/I hold194/I _7350_/Q _6333_/A1 _7801_/Q _4049_/A1 VDD VSS
+ gf180mcu_fd_sc_mcu7t5v0__aoi222_1
XFILLER_83_144 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_25_712 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7806_ _7806_/D _7877_/RN _7809_/CLK _7806_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffsnq_1
XPHY_206 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_52_531 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_239 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_228 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_217 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
X_5998_ _6547_/A1 _6004_/A2 _5998_/B hold432/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_4949_ _4951_/B _4979_/A3 _5458_/C VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_2
X_7737_ _7737_/D _7923_/RN _7737_/CLK _7737_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
X_7668_ _7668_/D _7923_/RN _7791_/CLK _7668_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffsnq_1
XFILLER_149_69 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_138_658 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_123_6 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6619_ _7918_/Q _6621_/A2 _6620_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_152_105 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7599_ hold94/Z _7923_/RN _7599_/CLK hold92/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_4_605 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_165_499 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_79_428 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
Xoutput280 _7349_/Q pll_trim[18] VDD VSS gf180mcu_fd_sc_mcu7t5v0__buf_4
XFILLER_0_811 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_58_22 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_121_558 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_94_409 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
Xoutput291 _7367_/Q pll_trim[4] VDD VSS gf180mcu_fd_sc_mcu7t5v0__buf_4
XFILLER_87_461 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_59_152 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_90_615 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_90_626 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_28_561 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_43_531 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_90_53 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_15_288 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_169_783 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_168_282 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_156_444 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_117_809 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_128_179 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_171_425 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_109_382 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_99_73 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_7_487 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_124_341 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_99_84 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_151_160 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_140_812 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_3_682 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_715 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_704 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_124_396 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_726 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_737 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_748 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_759 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_120_591 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_65_144 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6970_ _7862_/Q _7200_/B1 _7205_/B1 _7740_/Q _6971_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_5921_ hold500/Z _5936_/A2 hold501/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_34_531 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_46_380 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_5852_ _5852_/A1 hold5/Z _5853_/S VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_110_19 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_179_558 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_167_709 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5783_ _5104_/B _5783_/A2 _5783_/B _5783_/C _5784_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi211_1
X_4803_ _7488_/Q _4809_/S _4804_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_4734_ _7450_/Q hold50/Z _4741_/S hold51/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_7522_ _7522_/D _7961_/RN _7572_/CLK _7522_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_147_444 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_119_17 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_108_809 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_7453_ _7453_/D _7853_/RN _7461_/CLK _7453_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
X_4665_ _4685_/A1 hold558/Z _4665_/B hold559/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_134_105 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_147_499 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xhold900 hold900/I _7356_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
X_4596_ _6539_/A1 _4598_/A2 _4596_/B _7401_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
Xhold922 _7693_/Q hold922/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
Xhold911 _7701_/Q hold911/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
X_6404_ hold873/Z _6417_/A2 _6405_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_7384_ _7384_/D _7875_/RN _7790_/CLK _7384_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_162_469 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
Xhold955 _7412_/Q _4378_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
X_6335_ _6539_/A1 _6349_/A2 _6335_/B _7798_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
Xhold933 _7554_/Q _3635_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
Xhold944 _7555_/Q _3634_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
Xhold966 hold30/I hold966/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
XFILLER_0_107 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_88_247 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_8005_ _8005_/I _8005_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_6266_ hold845/Z _6281_/A2 _6267_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_5217_ _5392_/A1 _5254_/A3 _5218_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_6197_ hold638/Z _6208_/A2 hold639/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_69_472 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_69_461 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5148_ _5369_/B _5040_/B _5552_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_111_580 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_28_25 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_57_645 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5079_ _5087_/B _5456_/A2 _5079_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_84_486 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_84_475 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_56_188 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_12_203 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_44_46 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_40_534 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_12_247 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_166_753 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_100_96 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_60_34 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_181_712 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_176_34 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_180_211 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_165_296 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_153_425 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_114_2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_153_469 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_140_108 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_122_812 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_663 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_85_42 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_47_144 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_141_70 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_16_531 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_16_575 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_16_597 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_129_411 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_129_455 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_129_499 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_116_105 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xhold207 _7643_/Q hold207/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
X_4450_ _4487_/A1 _6539_/A1 _4450_/B _7347_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
Xhold218 hold218/I _7753_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
X_4381_ _7965_/Q _7964_/Q _4327_/S _3738_/Z _4383_/A1 _7414_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai32_1
Xhold229 _7987_/I hold229/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
XFILLER_7_295 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6120_ hold701/Z _6123_/A2 hold702/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_98_534 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_534 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_523 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_512 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_501 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_6051_ _4476_/I _6055_/A2 _6051_/B hold226/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
XTAP_545 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_556 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_567 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_5002_ _3723_/I _5662_/A1 _5643_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_4
XTAP_578 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_589 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_93_283 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6953_ _6953_/A1 _6953_/A2 _6955_/A4 _7202_/B1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor3_4
X_5904_ hold367/Z _5919_/A2 hold368/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_6884_ _7372_/Q _6644_/Z _6884_/B1 _7522_/Q _6886_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_5835_ _7566_/Q _5840_/A2 _5836_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_22_534 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_179_388 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5766_ _5766_/A1 _5766_/A2 _5766_/A3 _5767_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor3_1
XFILLER_163_712 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4717_ hold8/Z _3819_/Z _4717_/B _4718_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_5697_ _5419_/B _5697_/A2 _5697_/A3 _5697_/A4 _5698_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor4_1
X_7505_ _7505_/D _7961_/RN _7505_/CLK _7505_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
X_4648_ _4652_/A1 _4648_/A2 _4648_/B hold762/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_135_425 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_107_105 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_7436_ _7436_/D _7923_/RN _7599_/CLK _7436_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_30_37 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_163_778 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
Xhold730 _7455_/Q hold730/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
XFILLER_146_37 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_135_469 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_122_108 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_116_672 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_104_812 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7367_ _7367_/D _7875_/RN _7874_/CLK _7367_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffsnq_1
X_4579_ _4579_/A1 _6537_/A2 _4583_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
Xhold752 _7507_/Q hold752/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
Xhold763 _7409_/Q hold763/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
Xhold741 _7383_/Q hold741/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
X_7298_ _7901_/RN _4334_/Z _7298_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__and2_1
X_6318_ _6539_/A1 _6332_/A2 _6318_/B _7790_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
Xhold796 _7538_/Q hold796/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
Xhold774 _7373_/Q hold774/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
Xhold785 _7886_/Q hold785/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
XFILLER_89_567 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_77_729 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6249_ hold790/Z _6264_/A2 _6250_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_39_68 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_29_144 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_57_442 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_176_4 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_84_250 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xclkbuf_leaf_61_csclk clkbuf_3_3__f_csclk/Z _7820_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_72_434 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_41_810 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_111_73 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_71_22 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_13_512 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_13_567 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xclkbuf_leaf_76_csclk _7528_/CLK _7876_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_40_331 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_166_550 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_154_701 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_139_775 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_126_447 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_181_597 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_154_789 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_141_428 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_113_108 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_4_276 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_122_620 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
Xclkbuf_leaf_14_csclk _7873_/CLK _7864_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_121_141 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_110_804 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_121_163 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_95_548 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xclkbuf_leaf_29_csclk _7873_/CLK _7851_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
Xhold90 hold90/I hold90/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
XFILLER_48_486 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_75_283 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3950_ _7626_/Q _5954_/A1 _6073_/A1 _7682_/Q _4176_/C _3953_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi221_2
X_3881_ _3783_/Z _3925_/A2 hold75/Z _3963_/A4 _3881_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__or4_2
X_5620_ _5681_/A1 _5722_/A1 _5620_/B _5632_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_157_561 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5551_ _5644_/A2 _5739_/A2 _5551_/A3 _5557_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_77_2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_145_712 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_117_425 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4502_ hold233/Z _4504_/A2 _4502_/B hold472/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_172_531 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_145_778 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5482_ _5648_/A1 _5608_/B _5648_/B2 _5482_/B2 _5644_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_7221_ _7221_/A1 _7228_/S _7221_/B _7943_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_6_61 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_172_575 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_132_417 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_104_108 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_4433_ _7587_/Q input39/Z _4433_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__and2_1
X_4364_ _5224_/A3 _5224_/A4 _5302_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_7152_ _7797_/Q _7190_/A2 _7196_/A2 _7893_/Q _7153_/A4 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_4295_ _7339_/Q _4294_/Z _4308_/S VDD VSS gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_140_450 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_7083_ _7936_/Q _7133_/S _7109_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_59_718 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6103_ hold705/Z _6106_/A2 hold706/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_112_163 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6034_ _4476_/I _6038_/A2 _6034_/B hold356/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
XTAP_375 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_112_196 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_100_347 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_397 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_386 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_66_272 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_66_250 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2209 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_7985_ _7985_/I _7985_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_27_637 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_54_445 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1519 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1508 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_82_798 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_6936_ _6936_/A1 _6936_/A2 _6954_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_2
XPHY_26 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_15 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_37 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_26_169 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_54_478 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_168_804 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_81_286 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_48 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_59 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_179_174 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_179_141 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_22_331 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_6867_ _6867_/A1 _6867_/A2 _6867_/A3 _6867_/A4 _6867_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__and4_1
X_6798_ _7843_/Q _6894_/A2 _6659_/Z _7625_/Q _6890_/B1 _7851_/Q _6799_/A4 VDD VSS
+ gf180mcu_fd_sc_mcu7t5v0__aoi222_1
XFILLER_10_504 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5818_ hold772/Z _5827_/A2 _5819_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_50_673 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5749_ _5749_/A1 _5749_/A2 _5749_/A3 _5749_/A4 _5754_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand4_1
XFILLER_182_317 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_136_756 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_151_704 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_123_428 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_123_406 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7419_ _7419_/D _7853_/RN _7419_/CLK _7993_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
Xhold560 _7436_/Q hold560/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
XFILLER_151_759 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_150_247 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xhold571 _7726_/Q hold571/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
XFILLER_1_224 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_2_747 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xhold593 _7888_/Q hold593/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
Xhold582 _7622_/Q hold582/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
XFILLER_103_163 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_77_515 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_181_2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_85_570 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_57_272 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_57_283 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_82_32 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_60_459 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_158_325 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_15_70 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_9_357 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_127_712 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_126_211 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4080_ _4080_/A1 _4080_/A2 _4080_/A3 _4107_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_36_401 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_48_250 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_48_294 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_36_478 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4982_ _3722_/I _5006_/B _5254_/A2 _5662_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand3_4
X_7770_ _7770_/D _7901_/RN _7866_/CLK _7770_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_63_286 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_17_692 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_6721_ _7694_/Q _6881_/B1 _6721_/B _6721_/C _6729_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi211_1
X_3933_ _7876_/Q _6486_/A1 _6022_/A1 _7658_/Q _3936_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_23_139 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_32_640 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3864_ _3801_/Z _3864_/A2 hold81/Z _3864_/A4 hold149/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand4_4
X_6652_ _7838_/Q _6894_/A2 _6887_/B1 _7676_/Q _6683_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_5603_ _5603_/A1 _4993_/B _5753_/A2 _5798_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor3_1
X_3795_ _3810_/S hold579/Z _3795_/B _3963_/A4 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi21_4
XFILLER_118_734 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_6583_ _7908_/Q _6586_/A1 _6586_/B _6584_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand3_1
X_5534_ _5752_/C _5534_/A2 _5534_/A3 _5644_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor3_1
XFILLER_172_350 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5465_ _5465_/A1 _5803_/A1 _5772_/A3 _5799_/A1 _5472_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand4_1
X_4416_ _3810_/S _4416_/A2 _5903_/A2 _4416_/B2 _4416_/ZN VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai22_1
XFILLER_160_534 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_105_428 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7204_ _7400_/Q _7204_/A2 _7204_/B1 _7390_/Q _7208_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_132_269 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_132_247 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5396_ _5585_/A1 _5672_/A2 _5624_/B _5759_/A1 _5586_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_7135_ _7001_/C _7937_/Q _7161_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_141_792 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4347_ _7903_/Q _4347_/A2 _4360_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_7066_ _7898_/Q _7197_/A2 _7196_/A2 _7890_/Q _7196_/B1 _7640_/Q _7068_/A3 VDD VSS
+ gf180mcu_fd_sc_mcu7t5v0__aoi222_1
X_4278_ _7878_/Q _6503_/A1 _4719_/A1 input61/Z _4279_/A4 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_86_389 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_67_570 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6017_ _6549_/A1 _6021_/A2 _6017_/B _7649_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
XTAP_2006 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_27_412 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_27_434 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_39_283 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_39_294 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_55_732 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2039 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2017 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2028 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1305 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_70_702 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_36_69 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7968_ _7968_/D _7321_/Z _7972_/CLK hold62/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
Xclkbuf_1_0__f_wbbd_sck clkbuf_0_wbbd_sck/Z _3666__1/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XTAP_1338 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1327 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1316 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_14_128 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_55_798 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_153_6 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7899_ _7899_/D _7901_/RN _7899_/CLK _7899_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XTAP_1349 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_6919_ _7914_/Q _7913_/Q _6950_/A1 _6941_/A2 _7195_/B1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor4_4
XFILLER_167_144 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_128_509 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_182_103 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_109_712 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_108_200 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_182_136 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_136_531 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_108_211 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_10_378 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_136_575 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
Xhold390 _7812_/Q hold390/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
XFILLER_7_2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_151_589 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_77_312 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_77_87 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_93_42 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_73_540 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_18_445 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_93_97 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_45_286 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1861 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1850 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_61_768 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_159_645 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_159_623 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_1894 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1883 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1872 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_60_267 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_14_662 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_154_350 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_142_534 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5250_ _5779_/A1 _5425_/B _5783_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_114_247 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_69_802 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4201_ _4201_/A1 _4201_/A2 _4202_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_5181_ _5648_/A1 _5066_/Z _5608_/B _5186_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_4132_ _4075_/B _3847_/Z _5812_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_2
XFILLER_3_73 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_96_676 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_95_153 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_4063_ _4063_/A1 _4063_/A2 _4063_/A3 _4063_/A4 _4068_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand4_1
XFILLER_68_389 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_49_570 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_56_518 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_37_721 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_37_776 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_7822_ _7822_/D _7875_/RN _7822_/CLK _7822_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffsnq_1
XFILLER_37_798 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_51_212 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7753_ _7753_/D _7877_/RN _7755_/CLK _7753_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
X_4965_ _5797_/B _5363_/A2 _4965_/B _4969_/C VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi21_2
X_3916_ _3916_/A1 _3916_/A2 _3916_/A3 _3916_/A4 _3917_/A4 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand4_1
XFILLER_51_278 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6704_ _7749_/Q _6644_/Z _6884_/B1 _7685_/Q _6705_/A4 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_149_144 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7684_ _7684_/D _7923_/RN _7736_/CLK _7684_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffsnq_1
X_4896_ hold796/Z _4897_/A2 hold797/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_3847_ hold26/Z hold41/Z hold75/Z hold71/Z _3847_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__or4_4
XFILLER_20_676 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6635_ _6878_/A2 _6664_/A2 _6661_/A3 _6883_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor3_4
X_3778_ _3778_/I _7964_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_6566_ _6567_/A1 _6561_/Z _6567_/B1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_180_629 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_145_361 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5517_ _5517_/A1 _5642_/A3 _5517_/A3 _5517_/A4 _5518_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand4_1
XFILLER_105_225 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6497_ hold709/Z _6502_/A2 _6498_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_154_37 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5448_ _5448_/A1 _5777_/A2 _5448_/B _5461_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_133_567 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_133_545 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_105_236 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5379_ _5714_/A1 _5689_/A1 _5543_/C _5452_/C _5380_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi211_2
XFILLER_59_312 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7118_ _7698_/Q _7194_/A2 _7194_/B1 _7666_/Q _7194_/C1 _7812_/Q _7121_/A2 VDD VSS
+ gf180mcu_fd_sc_mcu7t5v0__aoi222_1
X_7049_ _7777_/Q _7200_/A2 _7193_/B1 _7631_/Q _7053_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_170_25 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_28_743 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_47_79 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_27_231 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_103_63 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_1113 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1102 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_27_286 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_82_392 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1146 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1124 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1135 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_63_34 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_15_437 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_144_2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1179 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1168 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1157 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_63_89 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_11_621 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_23_481 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_155_114 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_7_647 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_171_629 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_10_197 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_136_394 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_124_534 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_109_586 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_6_179 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_2_330 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_908 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_112_729 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_97_418 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_919 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_111_239 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_78_676 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_77_164 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_80_318 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_19_798 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_33_212 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2370 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_179_729 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_179_707 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_73_392 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_61_554 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2392 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2381 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_159_453 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4750_ hold729/Z _4750_/I1 _4753_/S _7463_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XTAP_1691 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1680 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_174_412 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4681_ _4685_/A1 hold521/Z _4681_/B hold522/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_146_103 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_119_306 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3701_ _7695_/Q _3701_/ZN VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_3632_ _3632_/I _3760_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_6420_ _6539_/A1 _6434_/A2 _6420_/B _7838_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_161_106 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6351_ hold489/Z _6366_/A2 _6352_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_5302_ _5302_/A1 _5011_/B _5302_/A3 _5319_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand3_2
XFILLER_115_523 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_115_512 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_170_662 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_115_567 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6282_ _6282_/A1 hold5/Z _6298_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_4
XFILLER_88_407 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_170_684 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5233_ _5254_/A2 _5616_/A1 _5365_/B1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_2
XFILLER_88_418 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5164_ _4993_/C _5452_/C _5543_/C _5559_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor3_2
XFILLER_110_250 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_84_602 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4115_ hold82/Z _4155_/A2 _7285_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_5095_ _5669_/A1 _5658_/B _5608_/B _4996_/Z _5095_/C _5098_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi221_1
XFILLER_96_495 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_68_197 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4046_ _4046_/A1 _4046_/A2 _4046_/A3 _4046_/A4 _4058_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand4_1
XFILLER_140_39 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_83_167 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7805_ _7805_/D _7853_/RN _7805_/CLK _7805_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XPHY_207 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_64_392 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_229 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_218 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
X_5997_ hold430/Z _6004_/A2 hold431/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_25_779 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_52_565 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4948_ _4944_/Z _4955_/A2 _5741_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_4
X_7736_ _7736_/D _7923_/RN _7736_/CLK _7736_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
X_7667_ _7667_/D _7853_/RN _7726_/CLK _7667_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
X_4879_ hold735/Z _4882_/A2 hold736/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_177_283 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_165_423 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6618_ _7435_/Q _7433_/Q _6618_/A3 _6618_/B _6621_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai31_1
X_7598_ _7598_/D _7853_/RN _7818_/CLK _7598_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_152_117 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_106_534 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6549_ _6549_/A1 _6553_/A2 _6549_/B _7899_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
Xoutput270 _7565_/Q pll_sel[2] VDD VSS gf180mcu_fd_sc_mcu7t5v0__buf_4
Xoutput292 _7368_/Q pll_trim[5] VDD VSS gf180mcu_fd_sc_mcu7t5v0__buf_4
Xoutput281 _7350_/Q pll_trim[19] VDD VSS gf180mcu_fd_sc_mcu7t5v0__buf_4
XFILLER_58_34 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_101_283 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_90_605 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_75_668 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_74_33 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_62_318 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_15_234 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_15_223 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_15_212 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_130_83 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_90_43 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_168_261 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_168_250 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_156_401 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_128_103 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_129_637 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_23_70 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_156_456 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_139_70 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_143_139 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_125_810 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_109_361 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_7_499 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_7_477 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_99_96 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_152_684 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_152_673 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_151_150 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_97_215 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_716 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_705 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_112_548 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_31_6 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_727 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_738 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_749 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_66_602 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_19_540 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_81_638 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5920_ _5920_/A1 _7285_/A2 _5936_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_4
XFILLER_0_85 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_46_392 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5851_ hold47/Z _5851_/A2 _5851_/B hold481/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_34_554 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5782_ _5782_/A1 _5782_/A2 _5782_/A3 _5795_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_21_215 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_4802_ _7221_/A1 _4809_/S _4802_/B _7487_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_4733_ _3830_/Z _4742_/A2 _4741_/S VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_4
X_7521_ _7521_/D _7961_/RN _7876_/CLK _7521_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_159_283 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7452_ hold35/Z _7853_/RN _7461_/CLK hold34/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
X_4664_ hold557/Z _3879_/Z _4664_/B hold558/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_119_169 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6403_ _6539_/A1 _6417_/A2 _6403_/B _7830_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_135_629 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_134_128 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4595_ hold756/Z _4598_/A2 _4596_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
Xhold901 _7767_/Q hold901/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
X_7383_ _7383_/D _7875_/RN _7790_/CLK _7383_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
Xhold912 hold912/I _6128_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
Xhold934 hold49/I hold934/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
X_6334_ hold784/Z _6349_/A2 _6335_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
Xhold945 hold945/I _7555_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
Xhold923 hold923/I _6111_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
Xhold967 hold11/I hold967/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
Xhold956 _7978_/Q _3736_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
XFILLER_131_802 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6265_ _6265_/A1 hold5/Z _6281_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_4
X_5216_ _5200_/B _3727_/I _5369_/B _5421_/B1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand3_2
XFILLER_142_194 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_8004_ _8004_/I _8004_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_97_760 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6196_ _4454_/Z _6208_/A2 _6196_/B hold918/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_5147_ _5528_/A2 _5020_/Z _5153_/C VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_2
XFILLER_130_389 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_111_570 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_28_37 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5078_ _3722_/I _5392_/A1 _5456_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_2
XFILLER_84_465 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_72_605 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4029_ input48/Z _4275_/A2 _5920_/A1 _7608_/Q _4030_/A4 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_44_318 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_37_392 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_52_362 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_100_31 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_9_709 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7719_ hold91/Z _7853_/RN _7722_/CLK _7719_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_165_286 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_153_415 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_107_810 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_109_73 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_107_2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_106_342 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_134_662 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_134_673 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_133_150 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_79_215 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_4_469 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_48_602 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_87_270 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_85_54 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_36_808 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_63_638 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_28_392 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_169_570 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_129_401 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_157_732 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_11_292 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_7_241 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_171_212 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_157_798 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xhold208 hold208/I _6004_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
Xhold219 _7601_/Q hold219/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
X_4380_ _4292_/B _4380_/A2 _4380_/B _7415_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_112_323 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_524 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_513 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_502 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_6050_ hold225/Z _6055_/A2 _6051_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_140_676 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_546 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_535 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_557 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_39_602 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_112_389 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5001_ _5600_/A1 _5363_/A2 _5663_/A1 _5585_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor3_2
XTAP_568 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_579 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_22_2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_38_134 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_26_307 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_54_605 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_121_19 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_81_424 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6952_ _6953_/A1 _6599_/Z _6955_/A4 _7204_/B1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor3_4
X_5903_ _5903_/A1 _5903_/A2 _7285_/A2 _5919_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand3_4
X_6883_ _7406_/Q _6883_/A2 _6883_/B1 _7398_/Q _6886_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_61_170 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5834_ _4460_/Z _5840_/A2 _5834_/B _7565_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_148_743 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5765_ _5765_/A1 _5765_/A2 _5765_/A3 _5766_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_175_540 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4716_ _3819_/Z hold2/Z _4717_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_148_754 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_147_242 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5696_ _5686_/Z _5696_/A2 _5695_/Z _5697_/A4 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand3_1
X_7504_ _7504_/D _7938_/RN _7638_/CLK _7504_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
X_4647_ _7456_/Q _3830_/Z _4647_/B _4648_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_147_286 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_107_128 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7435_ _7435_/D _7938_/RN _7940_/CLK _7435_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_2
Xhold720 _7827_/Q hold720/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
X_7366_ _7366_/D _7875_/RN _7875_/CLK _7366_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffsnq_1
XFILLER_162_267 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
Xhold731 _7380_/Q hold731/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
XFILLER_116_662 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_116_651 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6317_ hold794/Z _6332_/A2 _6318_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
Xhold742 _7368_/Q hold742/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
Xhold764 _7371_/Q hold764/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
Xhold753 _7389_/Q hold753/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
X_4578_ _4454_/Z _4578_/A2 _4578_/B _7394_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_7297_ _7877_/RN _4334_/Z _7297_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__and2_1
Xhold786 _7774_/Q hold786/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
Xhold797 hold797/I _4897_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
Xhold775 _7556_/Q hold775/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
XFILLER_1_428 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_39_14 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_130_131 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_130_142 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6248_ _6248_/A1 hold5/Z _6264_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_4
XFILLER_162_37 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_162_59 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6179_ _4454_/Z _6191_/A2 _6179_/B _7725_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_18_808 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_55_35 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_45_638 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_158_529 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_158_507 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_40_321 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_40_387 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_139_765 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_153_212 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_5_712 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_181_587 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_107_651 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_122_632 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_106_172 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_136_93 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_122_676 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_95_505 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_121_153 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_96_64 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_461 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_96_97 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
Xhold91 hold91/I hold91/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
Xhold80 hold80/I hold80/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
XFILLER_36_605 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_90_254 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_44_693 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_71_490 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3880_ hold609/Z hold42/Z _6469_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_4
XFILLER_176_337 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_31_354 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_129_231 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5550_ _5179_/B _5672_/A2 _5550_/B _5550_/C _5551_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XFILLER_172_510 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_172_521 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_157_584 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_129_286 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_5481_ _5658_/B _5179_/B _5757_/B _5765_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_4501_ hold470/Z _4504_/A2 hold471/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_7220_ _7943_/Q _7228_/S _7221_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_8_594 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_4432_ _7586_/Q input70/Z _4432_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_99_800 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_172_598 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4363_ _5302_/A1 _5195_/B _4906_/S VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_2
XFILLER_153_790 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_116_19 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_7151_ _7691_/Q _7189_/B1 _7189_/C1 _7659_/Q _7153_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_98_321 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4294_ hold87/I _7337_/Q _7336_/Q _4294_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__and3_1
X_6102_ _4476_/I _6106_/A2 _6102_/B hold334/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_112_120 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7082_ _7133_/S _7082_/A2 _7082_/B _7935_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_59_708 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6033_ hold355/Z _6038_/A2 _6034_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_376 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_398 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_387 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_7984_ _7984_/I _7984_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_1509 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_82_788 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6935_ _6941_/A2 _6935_/A2 _7190_/C1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_4
XPHY_27 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_16 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_38 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_23_800 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_49 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_22_321 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6866_ _7371_/Q _6644_/Z _6665_/Z _7537_/Q _6891_/C1 _7393_/Q _6867_/A4 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi222_1
X_6797_ _7795_/Q _6893_/A2 _6893_/B1 _7771_/Q _6893_/C1 _7633_/Q _6799_/A3 VDD VSS
+ gf180mcu_fd_sc_mcu7t5v0__aoi222_1
X_5817_ _5817_/A1 _6537_/A2 _5827_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_2
XFILLER_148_540 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5748_ _5748_/A1 _5748_/A2 _5777_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__or2_1
X_5679_ _5679_/A1 _5679_/A2 _5698_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_135_212 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_151_716 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7418_ _7418_/D _7853_/RN _7419_/CLK _7992_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
Xhold561 hold561/I _4690_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
Xhold572 _7992_/I hold572/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
Xhold550 _7704_/Q hold550/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
X_7349_ _7349_/D _7961_/RN _7505_/CLK _7349_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffsnq_1
XFILLER_89_354 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xhold594 hold594/I _6526_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
Xhold583 _7646_/Q hold583/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
XFILLER_131_473 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_104_676 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_77_527 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_66_34 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_58_741 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_18_605 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_58_763 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_174_2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_85_593 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_122_62 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_72_254 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_122_84 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_13_310 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_41_641 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_13_376 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_13_365 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_13_354 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_40_140 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_173_318 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_166_392 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_5_520 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_31_70 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_147_70 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_127_779 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_147_81 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_141_237 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_141_215 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_110_602 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_68_538 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_95_357 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_68_549 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_110_668 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_49_763 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_64_744 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4981_ _5309_/A1 _5709_/A1 _5777_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_4
XFILLER_17_682 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6720_ _6720_/A1 _6720_/A2 _6720_/A3 _6721_/C VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand3_1
X_3932_ _7730_/Q hold28/I _6124_/A1 _7706_/Q _6107_/A1 _7698_/Q _3936_/A1 VDD VSS
+ gf180mcu_fd_sc_mcu7t5v0__aoi222_1
X_3863_ _4075_/B _4151_/A2 _4249_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_4
XFILLER_32_685 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6651_ _7910_/Q _6664_/A2 _6661_/A3 _6887_/B1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor3_4
XFILLER_149_348 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5602_ _5602_/A1 _5602_/A2 _5797_/A2 _5602_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__or3_1
X_6582_ _7434_/Q _6585_/A2 _6590_/A1 _6587_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_164_318 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5533_ _5533_/A1 _5543_/B _5153_/C _5552_/A4 _5534_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor4_1
X_3794_ hold70/Z _3793_/Z _3810_/S hold71/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_4
XFILLER_118_724 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_145_521 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_117_212 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_172_340 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5464_ _5669_/B _5643_/A2 _5608_/B _4996_/Z _5799_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_1
Xclkbuf_leaf_60_csclk clkbuf_3_3__f_csclk/Z _7815_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
X_4415_ _3810_/S _4415_/A2 _4416_/B2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_5395_ _5669_/A1 _5783_/A2 _5685_/B _5292_/B _5703_/C _5398_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi221_1
X_7203_ _7404_/Q _7203_/A2 _7203_/B1 _7374_/Q _7208_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_99_641 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7134_ _7938_/Q _7133_/S _7161_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_4346_ _7435_/Q _4347_/A2 _6622_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_101_602 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_113_495 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_100_134 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_7065_ _7696_/Q _7194_/A2 _7194_/B1 _7664_/Q _7194_/C1 _7810_/Q _7068_/A2 VDD VSS
+ gf180mcu_fd_sc_mcu7t5v0__aoi222_1
Xclkbuf_leaf_75_csclk _7528_/CLK _7572_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
X_4277_ _7886_/Q _6520_/A1 _4527_/A1 _7373_/Q _4279_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_6016_ hold699/Z _6021_/A2 _6017_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_2007 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_100_189 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_36_37 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_2018 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2029 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_82_563 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_7967_ _7967_/D _7320_/Z _7972_/CLK hold30/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XTAP_1339 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1328 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1317 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1306 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_168_602 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6918_ _7914_/Q _7913_/Q _6936_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_2
X_7898_ _7898_/D _7900_/RN _7898_/CLK _7898_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_70_747 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_23_641 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_54_298 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_168_646 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_146_6 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6849_ _6849_/A1 _6767_/C _6849_/B1 _6849_/B2 _7433_/Q _6850_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi221_1
Xclkbuf_leaf_13_csclk clkbuf_leaf_9_csclk/I _7858_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_52_47 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_52_69 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_168_69 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_22_195 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_148_392 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xclkbuf_leaf_28_csclk _7873_/CLK _7773_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_124_738 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_123_226 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_123_215 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_151_579 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
Xhold380 hold380/I _7764_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
XFILLER_78_803 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_2_534 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_117_73 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_77_33 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
Xhold391 _7960_/Q hold391/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
XFILLER_77_357 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_46_744 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_45_276 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_1851 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1840 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_60_246 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1884 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1873 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1862 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_41_460 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_174_605 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_147_808 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1895 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_146_318 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_9_144 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_173_148 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_182_660 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_158_91 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4200_ _7807_/Q _6350_/A1 _4569_/A1 _7392_/Q _4812_/A1 _7495_/Q _4201_/A2 VDD VSS
+ gf180mcu_fd_sc_mcu7t5v0__aoi222_1
XFILLER_47_4 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5180_ _5648_/A1 _5774_/A1 _5752_/B1 _5066_/Z _5180_/C1 _5448_/A1 _5186_/A2 VDD VSS
+ gf180mcu_fd_sc_mcu7t5v0__aoi222_1
XFILLER_95_110 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4131_ _4141_/A1 _4217_/A2 _4893_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_4062_ hold98/I _6469_/A1 _4219_/A2 input14/Z _4063_/A4 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_110_498 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_64_530 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7821_ _7821_/D _7853_/RN _7821_/CLK _7821_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_36_276 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7752_ hold58/Z _7877_/RN _7752_/CLK hold57/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
X_4964_ _4965_/B _5363_/A2 _5774_/B2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_52_769 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_52_747 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3915_ _7683_/Q _6073_/A1 _6248_/A1 _7765_/Q _3916_/A4 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_6703_ _7661_/Q _6885_/A2 _6885_/B1 _7709_/Q _6705_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_177_454 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7683_ _7683_/D _7923_/RN _7698_/CLK _7683_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
X_4895_ hold47/Z _4897_/A2 _4895_/B hold395/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_165_638 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3846_ hold76/Z _4141_/A1 _6090_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_4
XFILLER_22_28 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6634_ _6634_/A1 _7906_/Q _6661_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_4
XFILLER_164_126 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_138_17 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3777_ input58/Z _3731_/Z _3777_/B1 _7964_/Q _3778_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_6565_ _6565_/A1 _6565_/A2 _6565_/B _7903_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_161_800 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_5516_ _5648_/A1 _5608_/B _5176_/B _5690_/A1 _5530_/B _5517_/A4 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi221_1
XFILLER_3_309 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6496_ _6547_/A1 _6502_/A2 _6496_/B hold535/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_173_682 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_160_321 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5447_ _5458_/C _5661_/A1 _5527_/A1 _5458_/B _5682_/A1 _5448_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai32_1
XFILLER_106_738 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_106_727 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_105_215 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_133_557 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_160_387 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5378_ _5585_/A1 _5708_/A2 _5378_/B _5378_/C _5733_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi211_2
XFILLER_99_460 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_87_600 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4329_ _4378_/B _4329_/A2 _7334_/Q _4330_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_7117_ _7852_/Q _7193_/A2 _7193_/B1 _7634_/Q _7193_/C1 _7730_/Q _7121_/A1 VDD VSS
+ gf180mcu_fd_sc_mcu7t5v0__aoi222_1
XFILLER_101_443 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7048_ _7048_/A1 _7048_/A2 _7048_/A3 _7048_/A4 _7054_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand4_1
XFILLER_59_357 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_59_368 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_170_37 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_86_176 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_28_733 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_90_809 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_27_221 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_1114 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1103 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_55_585 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_82_382 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1147 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1125 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1136 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1169 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1158 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_168_443 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_11_611 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_156_605 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_137_2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_128_307 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_10_132 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_149_690 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_10_176 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_7_637 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_171_619 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_109_565 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_151_354 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_88_32 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_2_375 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_909 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_120_741 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_92_102 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_92_179 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_80_308 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_18_276 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2371 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2360 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_34_747 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_2393 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2382 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_3700_ _7703_/Q _3700_/ZN VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XTAP_1692 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1681 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1670 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_14_460 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4680_ hold520/Z _3879_/Z _4680_/B hold521/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_147_638 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3631_ _7979_/Q _3735_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_143_800 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_6350_ _6350_/A1 hold5/Z _6366_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_4
XFILLER_155_693 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_5301_ _5301_/A1 _5303_/A4 _5301_/B _5359_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_52_2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_154_181 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_142_321 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6281_ _6553_/A1 _6281_/A2 _6281_/B _7773_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_5232_ _3722_/I _3723_/I _5006_/B _5006_/C _5303_/A4 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor4_4
X_5163_ _5319_/C _5692_/B _5645_/A1 _5501_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor3_1
XFILLER_142_398 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_96_463 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4114_ hold82/Z _3869_/I _4569_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_5094_ _5458_/B _5682_/A1 _5094_/B1 _5661_/A1 _5094_/C _5095_/C VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai221_1
XFILLER_68_187 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_84_669 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_84_658 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4045_ _7785_/Q _6299_/A1 hold28/I hold69/I _4249_/A2 input29/Z _4046_/A4 VDD VSS
+ gf180mcu_fd_sc_mcu7t5v0__aoi222_1
XFILLER_17_17 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_37_552 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_7804_ _7804_/D _7853_/RN _7851_/CLK _7804_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XPHY_219 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_208 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_12_408 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_24_246 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_24_268 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_25_769 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5996_ hold64/I _6004_/A2 _5996_/B hold181/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_4947_ _4943_/Z _4956_/A2 _4979_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_2
X_7735_ _7735_/D _7923_/RN _7735_/CLK _7735_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_33_780 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_138_605 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7666_ _7666_/D _7877_/RN _7812_/CLK _7666_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_20_441 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4878_ _4878_/A1 _6537_/A2 _4882_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_123_8 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3829_ hold609/I _3828_/I _4275_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_4
XFILLER_20_452 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_20_463 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_6617_ _7904_/Q _7905_/Q _6561_/Z _7435_/Q _6618_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai31_1
X_7597_ _7597_/D _7923_/RN _7597_/CLK _7597_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_165_37 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_152_129 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6548_ hold723/Z _6553_/A2 _6549_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_161_641 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6479_ _6547_/A1 _6485_/A2 _6479_/B hold436/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_160_140 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_133_354 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xoutput271 _7363_/Q pll_trim[0] VDD VSS gf180mcu_fd_sc_mcu7t5v0__buf_4
Xoutput260 _7571_/Q pll_bypass VDD VSS gf180mcu_fd_sc_mcu7t5v0__buf_4
XFILLER_133_387 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
Xoutput293 _7369_/Q pll_trim[6] VDD VSS gf180mcu_fd_sc_mcu7t5v0__buf_4
Xoutput282 _7364_/Q pll_trim[1] VDD VSS gf180mcu_fd_sc_mcu7t5v0__buf_4
XFILLER_59_154 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_101_273 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_87_496 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_74_124 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_28_541 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_28_530 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_74_179 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_16_747 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_31_706 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_90_55 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_90_33 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_31_728 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_129_627 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_90_88 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_90_66 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_11_496 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_7_434 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_137_682 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_99_64 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_136_192 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_124_321 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_98_717 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_706 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_155_70 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_97_227 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_717 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_728 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_739 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_78_463 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_78_441 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_120_582 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_66_636 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_38_316 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_93_499 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_80_105 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_65_157 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_80_116 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5850_ hold479/Z _5851_/A2 hold480/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_22_717 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_2190 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_5781_ _5565_/Z _5781_/A2 _5782_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_15_780 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4801_ _7487_/Q _4809_/S _4802_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_7520_ _7520_/D _7959_/RN _7545_/CLK _7520_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_4
X_4732_ _5903_/A2 _7285_/A2 _4742_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_2
X_7451_ hold14/Z _7853_/RN _7456_/CLK _7451_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
X_4663_ _3879_/Z _4460_/Z _4664_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_147_413 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_9_73 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_6402_ hold806/Z _6417_/A2 _6403_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_7382_ _7382_/D _7877_/RN _7849_/CLK _7382_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
Xhold902 _7564_/Q hold902/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
X_4594_ _4594_/A1 _6537_/A2 _4598_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
Xhold913 hold913/I _7701_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
Xhold935 hold935/I hold2/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
XFILLER_143_630 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_143_641 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6333_ _6333_/A1 hold5/Z _6349_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_4
Xhold946 _7553_/Q hold946/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
Xhold924 hold924/I _7693_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
Xhold957 hold1/I hold957/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
XFILLER_115_354 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6264_ _6553_/A1 _6264_/A2 _6264_/B hold254/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_5215_ _5200_/B _3727_/I _5421_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_8003_ _8003_/I _8003_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_6195_ hold916/Z _6208_/A2 hold917/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_5146_ _5643_/A2 _5752_/B1 _5186_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_97_783 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_69_496 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5077_ _5585_/A1 _5783_/A2 _5583_/C _5077_/C _5098_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi211_1
X_4028_ _7818_/Q _6367_/A1 _6265_/A1 _7770_/Q _4719_/A1 _8008_/I _4030_/A3 VDD VSS
+ gf180mcu_fd_sc_mcu7t5v0__aoi222_1
XFILLER_72_628 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_56_179 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_44_37 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_44_59 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_5979_ hold64/Z _5987_/A2 _5979_/B hold73/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_166_700 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_138_402 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7718_ _7718_/D _7853_/RN _7805_/CLK _7718_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffsnq_1
XFILLER_178_593 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_166_744 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_21_783 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
Xclkbuf_1_1__f__1040_ clkbuf_0__1040_/Z _7226_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
X_7649_ _7649_/D _7961_/RN _7649_/CLK _7649_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_60_58 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_109_52 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_106_321 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_109_96 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_109_85 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_69_34 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_79_227 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_69_89 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_121_357 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_95_709 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_632 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_125_73 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_85_44 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_48_636 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_87_282 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_47_146 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_62_105 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_75_499 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_62_116 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_16_522 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_71_672 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_70_171 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_43_363 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_176_508 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_34_70 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_7_231 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_172_747 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_125_641 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
Xhold209 hold209/I _7643_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
XFILLER_7_286 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_166_80 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_152_471 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_525 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_514 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_503 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_5000_ _5600_/A1 _5363_/A2 _5658_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_4
XTAP_547 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_536 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_558 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_79_783 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_569 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_15_2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_27_809 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_38_124 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_38_179 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6951_ _6955_/A4 _6951_/A2 _7188_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_4
XFILLER_81_458 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5902_ _6553_/A1 _5902_/A2 _5902_/B hold136/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_6882_ _7757_/Q _6882_/A2 _6882_/B1 _7495_/Q _6888_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_5833_ hold532/Z _5840_/A2 _5834_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_22_525 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_50_812 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_179_357 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5764_ _5579_/B _5764_/A2 _5744_/Z _5746_/Z _5805_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor4_2
X_7503_ _7503_/D _7503_/CLK _7503_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_4715_ hold131/Z _4718_/A1 hold132/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_148_766 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5695_ _5706_/A2 _5625_/Z _5725_/A2 _5691_/Z _5695_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__and4_1
X_4646_ _3830_/Z _4481_/I _4647_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_30_17 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7434_ _7434_/D _7938_/RN _7940_/CLK _7434_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_2
XFILLER_163_758 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
Xhold721 _7883_/Q hold721/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
Xhold710 _7796_/Q hold710/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
X_7365_ _7365_/D _7961_/RN _7567_/CLK _7365_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffsnq_1
X_4577_ hold861/Z _4578_/A2 _4578_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_162_257 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_150_408 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
Xhold732 _7779_/Q hold732/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
X_6316_ _6316_/A1 hold5/Z _6332_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_4
XFILLER_104_803 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xhold743 hold743/I _4517_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
Xhold754 _7399_/Q hold754/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
X_7296_ _7901_/RN _4334_/Z _7296_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__and2_1
Xhold787 _7862_/Q hold787/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
Xhold776 hold776/I _5814_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
Xhold765 _7580_/Q hold765/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
XFILLER_131_655 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_103_357 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_77_709 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xhold798 hold798/I _7538_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
X_6247_ _4454_/Z _6247_/A2 _6247_/B _7757_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_6178_ hold817/Z _6191_/A2 _6179_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_130_176 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_97_580 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_97_591 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5129_ _5705_/A2 _5179_/B _5657_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_85_731 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_69_282 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_85_775 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_44_105 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_57_499 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_111_31 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_111_53 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_25_374 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_41_812 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_111_97 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_138_210 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_166_552 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_166_530 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_139_755 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_154_703 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_154_747 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_126_438 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_107_641 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_181_566 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_134_460 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_106_140 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_5_779 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_4_267 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_122_611 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_121_132 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_106_195 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_121_176 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_96_54 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_29_70 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xhold92 hold92/I hold92/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
Xhold70 hold70/I hold70/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
Xhold81 hold81/I hold81/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
XFILLER_91_712 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_75_241 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_63_447 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_63_425 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_35_105 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_91_767 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_16_374 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_31_300 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_32_812 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_50_108 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_149_508 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5480_ _5538_/A1 _5026_/Z _5480_/A3 _5652_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_145_736 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_61_90 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4500_ _6549_/A1 _4504_/A2 _4500_/B hold747/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_4431_ input1/Z input36/Z _4431_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_132_408 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_99_812 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_153_780 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7150_ _7853_/Q _7193_/A2 _7189_/A2 _7715_/Q _7153_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_4362_ _6623_/B _4362_/A2 _7435_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_4293_ _4309_/S _4300_/C VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_6101_ hold332/Z _6106_/A2 hold333/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_7081_ _7935_/Q _7133_/S _7082_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_140_463 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_112_176 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_98_377 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6032_ _6547_/A1 _6038_/A2 _6032_/B _7656_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
XTAP_366 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_39_400 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_67_753 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_377 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_399 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_388 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_66_274 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_26_105 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_39_499 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7983_ _7983_/I _7983_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_6934_ _7912_/Q _7911_/Q _6941_/A2 _6908_/Z _7201_/B1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor4_4
XPHY_28 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_17 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_54_447 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_39 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_23_812 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_179_132 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_22_311 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6865_ _7756_/Q _6882_/A2 _6894_/C1 _7403_/Q _6865_/C _6867_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi221_1
X_6796_ _7763_/Q _6892_/A2 _6892_/B1 _7729_/Q _6799_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_5816_ _4454_/Z _5816_/A2 _5816_/B hold906/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_5747_ _5747_/A1 _5747_/A2 _5756_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_22_388 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5678_ _5678_/A1 _5064_/B _5678_/A3 _5679_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor3_1
XFILLER_136_747 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_108_427 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_7417_ _7417_/D _7853_/RN _7419_/CLK _7991_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
X_4629_ hold572/Z _4652_/A1 hold573/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_135_246 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
Xhold562 hold562/I _7436_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
Xhold540 hold540/I _5930_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
Xhold551 hold551/I _6134_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
X_7348_ _7348_/D _7961_/RN _7627_/CLK _7348_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffsnq_1
XFILLER_1_215 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_2_727 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
Xhold573 hold573/I _4632_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
X_7279_ _7279_/A1 _7279_/A2 _7279_/B _7517_/Q _7958_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi211_1
Xclkbuf_3_5__f_csclk clkbuf_0_csclk/Z _7422_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
Xhold595 hold595/I _7888_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
XFILLER_1_226 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xhold584 _7644_/Q hold584/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
XFILLER_106_53 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_103_176 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_77_539 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_73_712 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_45_425 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_167_2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_82_34 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_82_45 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_73_789 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_14_812 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_32_108 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_9_337 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_147_60 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_99_108 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_5_565 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_147_93 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_141_227 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_96_804 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_122_463 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_1_771 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
Xinput160 wb_rstn_i _7959_/RN VDD VSS gf180mcu_fd_sc_mcu7t5v0__buf_12
XFILLER_48_241 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_48_230 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_48_296 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_91_531 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4980_ _5741_/A1 _4993_/B _5735_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_4
XFILLER_51_428 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_3931_ _7674_/Q _6056_/A1 _5920_/A1 _7610_/Q _6367_/A1 _7820_/Q _3955_/A2 VDD VSS
+ gf180mcu_fd_sc_mcu7t5v0__aoi222_4
XFILLER_177_636 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3862_ hold26/Z hold41/Z hold75/Z hold71/Z _4151_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand4_4
XFILLER_31_141 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6650_ _6878_/A2 _6664_/A3 _6662_/A3 _6894_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor3_4
XFILLER_165_809 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5601_ _5783_/A2 _5668_/A2 _5668_/C _5612_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_82_2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_31_185 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6581_ _6586_/A1 _6581_/A2 _6663_/A4 _6586_/B _7907_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand4_1
XFILLER_176_179 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3793_ hold578/Z input58/Z _7414_/Q _3793_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_5532_ _5648_/A2 _5179_/B _5555_/B _5555_/C _5743_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XFILLER_118_747 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_117_224 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_11_19 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_145_566 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_118_769 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5463_ _5643_/A2 _5783_/A2 _5585_/B _5772_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_8_392 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xclkbuf_leaf_9_csclk clkbuf_leaf_9_csclk/I _7862_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_160_525 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_160_514 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5394_ _5394_/A1 _5709_/A2 _5394_/B _5415_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_4414_ _7919_/Q _7576_/Q _7580_/Q _4414_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_7202_ _7408_/Q _7202_/A2 _7202_/B1 _7398_/Q _7386_/Q _7202_/C2 _7208_/A1 VDD VSS
+ gf180mcu_fd_sc_mcu7t5v0__aoi222_1
X_7133_ _7133_/I0 _7937_/Q _7133_/S _7937_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_4345_ _7904_/Q _7905_/Q _4347_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_141_783 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_140_260 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7064_ hold59/I _7193_/A2 _7193_/B1 _7632_/Q _7193_/C1 _7728_/Q _7068_/A1 VDD VSS
+ gf180mcu_fd_sc_mcu7t5v0__aoi222_1
X_4276_ input52/Z _5886_/A1 _4888_/A1 _7535_/Q _4279_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_6015_ _6547_/A1 _6021_/A2 _6015_/B _7648_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_55_701 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_100_179 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_55_712 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2019 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2008 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_82_531 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7966_ _7966_/D _7319_/Z _7972_/CLK hold11/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XTAP_1329 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1318 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1307 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_14_108 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_42_406 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6917_ _6953_/A2 _6955_/A4 _6908_/Z _7207_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor3_4
X_7897_ _7897_/D _7900_/RN _7897_/CLK _7897_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffsnq_1
X_6848_ _6848_/A1 _6848_/A2 _6848_/A3 _6849_/B2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor3_1
XFILLER_22_130 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_52_37 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_168_669 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_168_37 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_139_6 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_23_697 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_23_686 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_52_59 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6779_ _7433_/Q _7924_/Q _6779_/B _6781_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_7_808 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_6_318 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_124_717 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_109_769 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_136_599 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_2_513 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_2_524 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
Xhold370 _7746_/Q hold370/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
Xhold381 _7985_/I hold381/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
XFILLER_123_238 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_117_41 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_89_130 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
Xhold392 _7666_/Q hold392/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
XFILLER_104_463 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_89_174 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_89_141 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_93_807 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_46_701 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_133_73 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_100_680 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_46_767 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_33_428 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_45_266 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1852 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1841 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1830 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_73_597 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1885 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1874 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1863 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_60_269 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_13_141 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1896 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_173_105 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_158_179 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_139_371 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_154_352 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_127_566 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_170_812 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_142_525 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_115_728 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_107_290 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_123_783 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_123_761 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_3_31 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4130_ hold82/Z _3881_/Z _4609_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_95_144 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4061_ input46/Z _4275_/A2 _5817_/A1 _7561_/Q _6282_/A1 _7777_/Q _4063_/A3 VDD VSS
+ gf180mcu_fd_sc_mcu7t5v0__aoi222_1
XFILLER_37_712 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7820_ _7820_/D _7923_/RN _7820_/CLK _7820_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
X_7751_ hold67/Z _7877_/RN _7755_/CLK hold66/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
X_4963_ _5069_/A2 _4930_/Z _4953_/Z _4963_/A4 _5363_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand4_4
X_3914_ _7731_/Q hold28/I _6384_/A1 _7829_/Q _3916_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_7682_ _7682_/D _7923_/RN _7820_/CLK _7682_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_32_450 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6702_ _6702_/A1 _6702_/A2 _6702_/A3 _6706_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_149_146 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_149_135 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4894_ hold393/Z _4897_/A2 hold394/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_20_601 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6633_ _7907_/Q _6633_/A2 _6665_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_165_628 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_164_105 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3845_ hold42/Z hold54/I hold43/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_4
XFILLER_22_18 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_177_499 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3776_ _7411_/Q _3730_/Z _4380_/A2 _3777_/B1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand3_1
X_6564_ _7435_/Q _6569_/A3 _6564_/B _7902_/Q _6565_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai211_1
X_5515_ _5179_/B _5672_/A2 _5550_/B _5517_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_6495_ hold533/Z _6502_/A2 hold534/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_161_812 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_133_503 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5446_ _5446_/A1 _5446_/A2 _5446_/A3 _5520_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_121_709 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_105_227 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_160_377 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5377_ _5378_/B _5711_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_59_303 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4328_ _7415_/Q _3734_/Z _4329_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_86_122 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7116_ _7116_/A1 _7116_/A2 _7116_/A3 _7116_/A4 _7130_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand4_1
X_7047_ _7655_/Q _7189_/C1 _7207_/B1 _7719_/Q _7048_/A4 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_4259_ _7660_/Q _6039_/A1 _5855_/A1 _7982_/I _4260_/A4 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_170_27 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_101_499 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_86_188 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_74_317 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_103_43 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1104 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_7949_ _7949_/D _7949_/CLK _7949_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_70_534 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1137 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1115 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1126 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_15_428 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_43_737 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1159 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_70_567 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1148 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_11_689 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_170_108 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_152_812 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_124_525 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_3_800 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_124_547 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_2_321 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_132_591 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_105_783 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_77_100 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_144_72 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_77_144 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_19_712 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_46_531 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_160_71 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_18_266 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_37_70 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_179_709 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2350 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2361 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_61_523 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2394 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2383 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2372 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1660 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_61_567 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_14_450 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1693 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1682 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1671 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_770 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_147_628 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
Xclkbuf_leaf_74_csclk _7528_/CLK _7650_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_159_499 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_146_105 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3630_ _7980_/Q _4424_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_161_108 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5300_ _5166_/C _5300_/A2 _5360_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_143_812 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6280_ hold273/Z _6281_/A2 _6281_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
Xclkbuf_leaf_89_csclk _7528_/CLK _7638_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_6_693 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_5_170 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5231_ _4915_/Z _5303_/A3 _5258_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_102_208 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_69_601 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_45_2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5162_ _5218_/B _5498_/B _5162_/B _5162_/C _5187_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai211_1
X_5093_ _5087_/C _4898_/Z _5424_/A1 _5094_/C VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand3_1
Xclkbuf_leaf_12_csclk clkbuf_leaf_9_csclk/I _7854_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
X_4113_ _3828_/I _4141_/A1 _4878_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_56_317 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4044_ _7687_/Q _6090_/A1 _6073_/A1 _7679_/Q _6141_/A1 hold84/I _4046_/A3 VDD VSS
+ gf180mcu_fd_sc_mcu7t5v0__aoi222_1
XFILLER_140_19 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
Xclkbuf_leaf_27_csclk _7873_/CLK _7829_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
X_7803_ _7803_/D _7853_/RN _7805_/CLK _7803_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_24_236 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_52_534 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_209 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
X_7734_ _7734_/D _7923_/RN _7734_/CLK _7734_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffsnq_1
XFILLER_24_258 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5995_ hold179/Z _6004_/A2 hold180/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_40_707 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_52_567 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4946_ _4946_/A1 _5230_/A1 _4917_/Z _5369_/B _4955_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai22_2
XFILLER_33_17 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_33_792 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_7665_ _7665_/D _7853_/RN _7726_/CLK _7665_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
X_4877_ _4454_/Z _4877_/A2 _4877_/B hold802/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_7596_ _7596_/D _7923_/RN _7600_/CLK _7596_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_165_425 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_137_105 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3828_ _3828_/I _4620_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_6616_ _7916_/Q _6611_/B _6616_/B _7916_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_137_138 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6547_ _6547_/A1 _6553_/A2 _6547_/B hold447/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_3759_ _4292_/B _3759_/A2 _7974_/Q _3760_/B2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_152_108 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_146_672 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_134_812 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_133_344 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_118_396 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_106_536 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6478_ hold434/Z _6485_/A2 hold435/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_5429_ _5624_/A1 _5648_/B2 _5685_/B _5614_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
Xoutput261 _7557_/Q pll_dco_ena VDD VSS gf180mcu_fd_sc_mcu7t5v0__buf_4
Xoutput250 _4435_/Z pad_flash_csb_oe VDD VSS gf180mcu_fd_sc_mcu7t5v0__buf_4
XFILLER_161_697 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
Xoutput272 _7357_/Q pll_trim[10] VDD VSS gf180mcu_fd_sc_mcu7t5v0__buf_4
Xoutput283 _7351_/Q pll_trim[20] VDD VSS gf180mcu_fd_sc_mcu7t5v0__buf_4
Xoutput294 _7370_/Q pll_trim[7] VDD VSS gf180mcu_fd_sc_mcu7t5v0__buf_4
XFILLER_59_144 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_114_31 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_74_57 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_16_737 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_90_12 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_43_567 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_169_720 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_130_85 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_70_386 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_169_775 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_156_403 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_90_78 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_11_442 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_128_105 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_171_428 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_143_119 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_125_812 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_109_363 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_151_141 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_3_641 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_707 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_718 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_31_8 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_729 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_39_807 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_171_70 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_93_456 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_93_445 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_74_692 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_87 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_34_534 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_46_372 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2180 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_61_353 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4800_ _7219_/A1 _4809_/S _4800_/B _7486_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
XTAP_2191 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_5780_ _5372_/Z _5780_/A2 _5780_/B _5781_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_175_712 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_159_241 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1490 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_4731_ _6549_/A1 _4731_/A2 _4731_/B _7449_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_7450_ hold51/Z _7853_/RN _7461_/CLK _7450_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_147_436 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_147_425 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4662_ _7983_/I _4685_/A1 _4665_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_30_751 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_174_244 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6401_ _6401_/A1 _6537_/A2 _6417_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_4
X_7381_ _7381_/D _7877_/RN _7381_/CLK _7381_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_134_108 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_128_672 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
Xhold903 _7871_/Q hold903/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
X_4593_ _4454_/Z _4593_/A2 _4593_/B _7400_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
Xhold936 hold21/I hold936/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
X_6332_ _6553_/A1 _6332_/A2 _6332_/B hold318/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_115_311 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
Xhold914 _7407_/Q hold914/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
Xhold925 _7791_/Q hold925/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
Xhold958 _3766_/Z _7972_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
X_6263_ hold252/Z _6264_/A2 hold253/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_89_707 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
Xhold947 _7550_/Q hold947/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
X_5214_ _5669_/A1 _5087_/B _5218_/C VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_88_239 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_8002_ _8002_/I _8002_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_6194_ hold47/Z _6208_/A2 _6194_/B hold674/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_5145_ _5643_/A2 _5608_/B _5739_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_111_561 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_111_550 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_97_795 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_96_250 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5076_ _5669_/B _4996_/Z _5465_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_84_445 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_4027_ _7744_/Q hold43/I _6248_/A1 _7762_/Q _4030_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_25_534 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_13_707 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_25_556 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_25_567 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5978_ _7631_/Q _5987_/A2 _5979_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_80_673 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4929_ _5195_/B _4914_/Z _5210_/A3 _4951_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor3_2
X_7717_ _7717_/D _7877_/RN _7747_/CLK _7717_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffsnq_1
XFILLER_100_55 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_20_250 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7648_ _7648_/D _7961_/RN _7960_/CLK _7648_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_60_37 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_176_37 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_176_15 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_165_244 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_181_737 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_176_59 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_153_428 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_153_406 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_107_812 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7579_ _7579_/D _7961_/RN _7624_/CLK _7579_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_180_247 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_109_64 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_134_664 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_122_804 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_106_388 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_688 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_699 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_75_445 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_75_456 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_141_73 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_16_534 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_157_712 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_156_211 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_156_200 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_129_425 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_157_778 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_12_795 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_11_283 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_8_744 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_116_108 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_8_788 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_125_620 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_109_160 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_124_130 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_515 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_504 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_140_656 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_112_347 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_548 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_537 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_526 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_79_795 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_78_250 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_559 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_120_380 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_94_743 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_66_445 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6950_ _6950_/A1 _6950_/A2 _6955_/A4 _7204_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor3_4
XFILLER_66_478 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_66_456 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_94_798 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_93_286 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5901_ hold134/Z _5902_/A2 hold135/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_6881_ _7530_/Q _6881_/A2 _6881_/B1 _7524_/Q _6888_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_62_673 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5832_ _4454_/Z _5840_/A2 _5832_/B _7564_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_22_504 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_22_515 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5763_ _5763_/A1 _5698_/B _5763_/A3 _5763_/A4 _5792_/B1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor4_2
XFILLER_14_19 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_4714_ _4718_/A1 hold530/Z _4714_/B hold531/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_7502_ _7502_/D _7503_/CLK _7502_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_5694_ _5424_/Z _5763_/A1 _5723_/A1 _5694_/A4 _5696_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor4_1
XFILLER_162_203 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4645_ hold761/Z _4652_/A1 _4648_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_135_428 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7433_ _7433_/D _7938_/RN _7940_/CLK _7433_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_4
XFILLER_162_247 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xhold711 _7610_/Q hold711/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
X_7364_ _7364_/D _7875_/RN _7875_/CLK _7364_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffsnq_1
X_4576_ _6539_/A1 _4578_/A2 _4576_/B _7393_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
Xhold700 _7449_/Q hold700/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
XFILLER_115_130 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_6315_ _6553_/A1 _6315_/A2 _6315_/B _7789_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
Xhold722 _7859_/Q hold722/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
Xhold755 _7504_/Q hold755/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
Xhold744 hold744/I _7368_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
Xhold733 _7352_/Q hold733/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
XFILLER_1_408 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7295_ _7877_/RN _4334_/Z _7295_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_115_152 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_89_515 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
Xhold777 hold777/I _7556_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
Xhold766 _7403_/Q hold766/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
Xhold788 _7894_/Q hold788/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
XFILLER_103_336 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
Xhold799 _7854_/Q hold799/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
X_6246_ hold815/Z _6247_/A2 _6247_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_6177_ hold47/Z _6191_/A2 _6177_/B _7724_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_97_570 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_85_721 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5128_ _5600_/A1 _5797_/B _5527_/A1 _5166_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor3_1
XFILLER_130_199 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_84_264 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_29_169 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5059_ _5195_/B _5016_/B _5692_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_4
XFILLER_85_798 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_57_489 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_72_459 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_111_65 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_40_301 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_139_712 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_21_570 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_40_389 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_138_266 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_112_2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_121_144 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_463 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_496 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_48_445 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xhold60 hold60/I hold60/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
Xhold71 hold71/I hold71/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
Xhold82 hold82/I hold82/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
XFILLER_91_702 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_29_82 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
Xhold93 hold93/I hold93/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
XFILLER_75_286 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_17_810 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_91_779 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_91_757 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_45_70 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_44_673 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_31_312 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_145_704 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_12_592 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_172_534 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_117_428 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4430_ _4396_/S input63/Z _4430_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_144_269 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_144_247 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_6_53 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_6100_ _6547_/A1 _6106_/A2 _6100_/B hold538/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_4361_ _7433_/Q _4361_/A2 _4361_/A3 _4362_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand3_1
X_4292_ _7414_/Q _4292_/A2 _4292_/B _4309_/S VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_4
XFILLER_112_122 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7080_ _7433_/Q _7934_/Q _7078_/Z _7080_/B2 _7082_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_112_155 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_98_389 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6031_ hold553/Z _6038_/A2 _6032_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_79_570 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_367 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_389 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_378 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_81_212 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7982_ _7982_/I _7982_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_26_128 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_54_426 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_54_437 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_6933_ _6941_/A2 _6951_/A2 _7193_/B1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_4
XPHY_18 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_29 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_54_459 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6864_ _6864_/A1 _6864_/A2 _6864_/A3 _6865_/C VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_179_144 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_90_790 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5815_ hold904/Z _5816_/A2 hold905/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_6795_ _7827_/Q _6891_/A2 _6891_/B1 _7673_/Q _6891_/C1 _7779_/Q _6799_/A1 VDD VSS
+ gf180mcu_fd_sc_mcu7t5v0__aoi222_1
XFILLER_50_676 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5746_ _5380_/I _5501_/Z _5524_/I _5746_/A4 _5746_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__or4_1
XFILLER_148_531 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_10_529 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_41_17 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_148_586 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_5677_ hold24/I _5520_/C _5677_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__and2_1
X_4628_ _4652_/A1 hold569/Z _4628_/B hold570/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_7416_ _7416_/D _7853_/RN _7419_/CLK _7990_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
Xhold530 hold530/I hold530/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
XFILLER_163_567 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_151_718 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_173_16 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
Xhold563 _7750_/Q hold563/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
XFILLER_150_206 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_144_770 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
Xhold541 hold541/I _7608_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
Xhold552 hold552/I _7704_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
X_7347_ _7347_/D _7961_/RN _7505_/CLK _7347_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffsnq_1
X_4559_ _4559_/A1 _6537_/A2 _4563_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_7278_ _7278_/A1 _7277_/B _7278_/B _7957_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi21_1
Xhold574 hold574/I _7418_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
Xhold585 _7760_/Q hold585/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
Xhold596 _7638_/Q hold596/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
X_6229_ hold831/Z hold6/Z _6230_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_103_144 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_77_529 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_890 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_57_286 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_45_459 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_82_57 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_26_673 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_15_73 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_13_367 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_40_131 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_139_564 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_139_553 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_154_534 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_126_269 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_126_258 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_126_247 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_68_529 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_68_518 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_95_337 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_282 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_1_783 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xinput150 wb_dat_i[2] _7252_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyb_1
Xinput161 wb_sel_i[0] _7236_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XFILLER_63_212 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_36_448 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3930_ _7884_/Q _6503_/A1 _5870_/A1 _3927_/Z _6005_/A1 _7650_/Q _3955_/A1 VDD VSS
+ gf180mcu_fd_sc_mcu7t5v0__aoi222_4
XFILLER_176_103 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3861_ hold27/Z _4141_/A1 hold28/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_4
XFILLER_32_676 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3792_ hold49/Z hold70/Z _3795_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__and2_1
X_5600_ _5600_/A1 _5797_/B _4993_/C _5458_/B _5600_/B2 _5668_/C VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai32_1
X_6580_ _7432_/Q _4352_/B _6586_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_2
XFILLER_173_810 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5531_ _5543_/B _5539_/A3 _5541_/A4 _5555_/C VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor3_2
XFILLER_75_2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5462_ _4969_/C _5604_/A2 _5658_/B _5608_/B _5462_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__or4_1
X_7201_ _7372_/Q _7201_/A2 _7201_/B1 _7508_/Q _7206_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_5393_ _5380_/I _5565_/A2 _5581_/C _5394_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__or3_1
X_4413_ _7917_/Q _7577_/Q _7580_/Q _4413_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_4344_ _4344_/I _7520_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_7132_ _7433_/Q _7132_/A2 _7132_/B _7133_/I0 VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_140_250 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_113_453 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7063_ _7063_/A1 _7063_/A2 _7063_/A3 _7063_/A4 _7078_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand4_1
XFILLER_98_175 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_86_315 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6014_ hold396/Z _6021_/A2 _6015_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_4275_ input43/Z _4275_/A2 _4549_/A1 _7383_/Q _4279_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_39_231 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_39_286 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_2009 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_94_392 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_82_543 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7965_ _7965_/D _7318_/Z _4415_/A2 _7965_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XTAP_1319 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1308 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_7896_ _7896_/D _7901_/RN _7896_/CLK _7896_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
X_6916_ _6950_/A1 _6941_/A2 _6908_/Z _7189_/B1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor3_4
XFILLER_70_749 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6847_ _6847_/A1 _6847_/A2 _6847_/A3 _6848_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_50_451 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_6778_ _7079_/A1 _6767_/C _6778_/B _7433_/Q _6779_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XFILLER_164_810 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5729_ _5791_/A2 _5761_/A2 _5762_/A4 _5730_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_50_495 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_136_534 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_108_247 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_108_269 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_117_31 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
Xhold371 _7804_/Q hold371/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
Xhold360 _7362_/Q hold360/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
Xhold382 hold382/I _4673_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
XFILLER_117_64 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_78_805 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_77_35 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xhold393 _7537_/Q hold393/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
XFILLER_131_283 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_131_272 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_131_294 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_92_318 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_93_34 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_85_381 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_18_459 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1842 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1831 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1820 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_159_615 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_158_103 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1875 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1864 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1853 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1897 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1886 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_14_676 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_155_810 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_139_361 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_9_168 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_154_342 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_182_684 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_182_695 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_127_578 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_122_250 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_96_602 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_96_635 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_95_112 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_95_123 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_4060_ _7615_/Q _5937_/A1 _6226_/A1 hold66/I _4063_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_76_392 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_37_735 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_64_554 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7750_ _7750_/D _7877_/RN _7755_/CLK _7750_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffsnq_1
X_4962_ _5369_/B _4943_/Z _5603_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_4
XFILLER_51_215 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3913_ _7715_/Q _6141_/A1 _6265_/A1 _7773_/Q _3916_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_7681_ _7681_/D _7853_/RN _7720_/CLK _7681_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
X_4893_ _4893_/A1 _7285_/A2 _4897_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_6701_ _7376_/Q _6882_/A2 _6880_/A2 _7815_/Q _6702_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_149_125 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_149_114 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3844_ _4212_/A2 _4075_/B _4488_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_4
X_6632_ _7910_/Q _6664_/A3 _6662_/A3 _6881_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor3_4
XFILLER_20_646 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_3775_ _7965_/Q _3738_/Z _4380_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_6563_ _6563_/I _6565_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_5514_ _5514_/A1 _5514_/A2 _5514_/A3 _5514_/A4 _5518_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand4_1
X_6494_ _6545_/A1 _6502_/A2 _6494_/B hold460/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_118_534 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_118_578 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_5445_ _5783_/B _5757_/B _5445_/A3 _5445_/A4 _5446_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor4_1
XFILLER_133_559 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_114_740 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5376_ _5371_/C _5392_/B2 _5376_/B _5378_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_7115_ _7690_/Q _7189_/B1 _7189_/C1 _7658_/Q _7115_/C _7116_/A4 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi221_1
XFILLER_160_389 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_141_570 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_4327_ _7964_/Q _7335_/Q _4327_/S _7335_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_113_283 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_101_423 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_101_412 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_86_112 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_101_445 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7046_ hold69/I _7193_/C1 _7196_/B1 _7639_/Q _7048_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_4258_ _7716_/Q hold90/I _4878_/A1 _7531_/Q _4260_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_103_33 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_67_392 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_27_212 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4189_ input72/Z _5903_/A1 _4232_/A2 input35/Z _4584_/A1 _7398_/Q _4203_/A3 VDD VSS
+ gf180mcu_fd_sc_mcu7t5v0__aoi222_2
XFILLER_82_340 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1105 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_55_554 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7948_ _7948_/D _7949_/CLK _7948_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_1138 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1116 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1127 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_151_6 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1149 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_7879_ _7879_/D _7900_/RN _7900_/CLK _7879_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffsnq_1
XFILLER_23_495 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_155_128 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_6_116 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_6_105 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_136_331 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_109_567 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_109_534 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_164_673 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_163_161 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_3_812 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_88_34 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_78_602 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_5_2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xhold190 _7659_/Q hold190/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
XFILLER_105_795 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_104_250 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_66_808 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_93_638 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_19_757 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_58_392 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xclkbuf_leaf_8_csclk clkbuf_leaf_9_csclk/I _7878_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_19_779 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2351 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2362 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2340 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_33_215 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_34_727 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2395 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2384 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2373 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1650 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1694 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1683 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1672 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1661 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_53_70 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_169_70 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_154_161 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_154_150 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_6_672 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_182_492 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5230_ _5230_/A1 _5054_/Z _5685_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_4
XFILLER_5_160 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_170_676 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_5161_ _3723_/I _5579_/B _5162_/C VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_142_389 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_123_570 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_38_2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_5092_ _5058_/Z _5456_/A2 _5114_/A3 _5776_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand3_2
XFILLER_84_605 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4112_ hold82/Z _3963_/Z _4614_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_111_798 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4043_ _7735_/Q _6192_/A1 _6124_/A1 _7703_/Q _6107_/A1 _7695_/Q _4046_/A2 VDD VSS
+ gf180mcu_fd_sc_mcu7t5v0__aoi222_1
XFILLER_68_156 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_49_392 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_80_811 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7802_ _7802_/D _7901_/RN _7858_/CLK _7802_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
X_5994_ _4460_/Z _6004_/A2 _5994_/B _7638_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_4945_ _4900_/Z _4915_/Z _4945_/B1 _5022_/B _4956_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_2
X_7733_ _7733_/D _7938_/RN _7733_/CLK _7733_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffsnq_1
XFILLER_52_546 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_178_743 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7664_ hold39/Z _7877_/RN _7849_/CLK _7664_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_149_29 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_60_590 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4876_ hold800/Z _4877_/A2 hold801/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_177_286 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_165_415 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_3827_ _3783_/Z _3925_/A2 hold75/Z hold71/Z _3828_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand4_4
X_7595_ _7595_/D _7900_/RN _7892_/CLK _8005_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
X_6615_ _7916_/Q _6586_/B _6611_/B _6616_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand3_1
X_3758_ _7975_/Q _3765_/A1 _3759_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_118_331 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6546_ hold445/Z _6553_/A2 hold446/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_180_407 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_165_17 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_146_662 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_173_492 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3689_ _7785_/Q _3689_/ZN VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_6477_ _6545_/A1 _6485_/A2 hold99/Z hold100/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_5428_ _5482_/B2 _5510_/A2 _5793_/B _5789_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi21_1
Xoutput262 _7558_/Q pll_div[0] VDD VSS gf180mcu_fd_sc_mcu7t5v0__buf_4
Xoutput251 _4423_/Z pad_flash_io0_do VDD VSS gf180mcu_fd_sc_mcu7t5v0__buf_4
Xoutput240 _7984_/Z mgmt_gpio_out[3] VDD VSS gf180mcu_fd_sc_mcu7t5v0__buf_4
X_5359_ _5359_/A1 _5359_/A2 _5636_/A1 _5359_/B _5360_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai31_1
Xoutput284 _7352_/Q pll_trim[21] VDD VSS gf180mcu_fd_sc_mcu7t5v0__buf_4
Xoutput273 _7358_/Q pll_trim[11] VDD VSS gf180mcu_fd_sc_mcu7t5v0__buf_4
Xoutput295 _7355_/Q pll_trim[8] VDD VSS gf180mcu_fd_sc_mcu7t5v0__buf_4
XFILLER_58_37 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7029_ _7933_/Q _7133_/S _7030_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_75_638 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_101_286 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_83_660 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_70_321 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_15_215 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_130_75 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_142_2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_70_398 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_7_414 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_23_73 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_156_448 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_139_73 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_128_139 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_7_436 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_7_425 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_152_676 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_155_83 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_155_94 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_105_570 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_2_174 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_708 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_719 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_2_185 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_78_487 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_66_605 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_38_318 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_66_638 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_171_82 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_65_159 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_19_554 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_80_118 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_73_170 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_77 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_19_576 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_2170 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2192 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2181 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1491 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1480 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_4730_ hold700/Z _4731_/A2 _4731_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_159_286 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4661_ _4685_/A1 _4661_/A2 _4661_/B hold619/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_9_97 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_175_779 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_159_297 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7380_ _7380_/D _7877_/RN _7877_/CLK _7380_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
X_6400_ _6553_/A1 _6400_/A2 _6400_/B hold262/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_162_418 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6331_ hold316/Z _6332_/A2 hold317/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
Xhold904 _7557_/Q hold904/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
X_4592_ hold838/Z _4593_/A2 _4593_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
Xhold937 _7956_/Q _3673_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
Xhold926 _7653_/Q hold926/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
Xhold915 _7815_/Q hold915/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
Xhold959 hold87/I hold959/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
X_6262_ hold233/Z _6264_/A2 _6262_/B hold380/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
Xhold948 _7549_/Q hold948/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
X_5213_ _4906_/Z _5373_/A3 _5373_/A4 _5405_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand3_4
X_8001_ hold95/I _8001_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_6193_ hold672/Z _6208_/A2 hold673/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_5144_ _5543_/C _5689_/A2 _5543_/B _5499_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor3_1
X_5075_ _5603_/A1 _4993_/B _5663_/A1 _5583_/C VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor3_2
XFILLER_57_638 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4026_ _7826_/Q _6384_/A1 hold150/I _7567_/Q _6537_/A1 _7898_/Q _4030_/A1 VDD VSS
+ gf180mcu_fd_sc_mcu7t5v0__aoi222_1
XFILLER_52_321 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5977_ _4460_/Z _5987_/A2 _5977_/B _7630_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_52_387 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4928_ _4914_/Z _5210_/A3 _5195_/B _5069_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_4
X_7716_ _7716_/D _7853_/RN _7726_/CLK _7716_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffsnq_1
XFILLER_100_45 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_40_538 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_165_212 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_100_89 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7647_ _7647_/D _7961_/RN _7960_/CLK hold78/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_165_234 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4859_ hold597/Z _4862_/A2 hold598/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_180_204 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_109_21 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_7578_ _7578_/D _7961_/RN _7624_/CLK _7578_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_119_695 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_118_183 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6529_ hold438/Z _6536_/A2 hold439/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_134_676 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_133_164 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_133_175 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_79_229 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_79_207 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_88_796 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_667 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_48_605 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xclkbuf_leaf_73_csclk _7528_/CLK _7961_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_28_384 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_71_641 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xclkbuf_leaf_88_csclk _7528_/CLK _7505_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_43_321 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_71_674 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_16_579 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_43_354 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xclkbuf_leaf_11_csclk clkbuf_leaf_9_csclk/I _7863_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_129_459 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_8_734 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_171_215 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_125_632 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xclkbuf_leaf_26_csclk _7422_/CLK _7872_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_124_142 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_109_194 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_140_602 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_516 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_505 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_549 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_538 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_527 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_120_392 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_78_273 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_39_638 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5900_ hold233/Z _5902_/A2 _5900_/B hold295/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_34_321 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_34_343 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6880_ _7961_/Q _6880_/A2 _6880_/B1 _7410_/Q _7477_/Q _6880_/C2 _6888_/A1 VDD VSS
+ gf180mcu_fd_sc_mcu7t5v0__aoi222_1
XFILLER_179_315 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5831_ hold902/Z _5840_/A2 _5832_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_5762_ _5776_/A1 _5778_/A1 _5762_/A3 _5762_/A4 _5763_/A4 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand4_1
XFILLER_34_387 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4713_ hold529/Z _3819_/Z _4713_/B hold530/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_7501_ _7501_/D _7503_/CLK _7501_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_147_212 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5693_ _5424_/Z _5694_/A4 _5762_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_175_565 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_163_716 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4644_ _4652_/A1 _4644_/A2 _4644_/B hold693/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_30_19 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7432_ _7432_/D _7961_/RN _7940_/CLK _7432_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffsnq_1
Xhold701 _7698_/Q hold701/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
Xhold712 _7682_/Q hold712/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
X_7363_ _7363_/D input75/Z _7567_/CLK _7363_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffsnq_1
X_4575_ hold771/Z _4578_/A2 _4576_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_7294_ _7901_/RN _4334_/Z _7294_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__and2_1
X_6314_ hold245/Z _6315_/A2 _6315_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
Xhold723 _7899_/Q hold723/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
Xhold734 _7472_/Q hold734/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
Xhold745 _7360_/Q hold745/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
XFILLER_170_270 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_116_676 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_89_527 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xhold756 _7401_/Q hold756/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
Xhold767 _7444_/Q hold767/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
Xhold778 _7405_/Q hold778/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
X_6245_ _6539_/A1 _6247_/A2 _6245_/B _7756_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
Xhold789 _7838_/Q hold789/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
XFILLER_162_29 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6176_ hold523/Z _6191_/A2 _6177_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_5127_ _5648_/A2 _5643_/A2 _5803_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_57_424 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5058_ _5195_/B _5016_/B _5058_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_29_159 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4009_ _7359_/Q _4488_/A1 _6124_/A1 _7704_/Q _4176_/C _4013_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi221_1
XFILLER_38_660 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_37_181 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_53_641 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_52_195 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_178_392 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_138_212 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_139_779 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_153_215 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_153_248 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_106_142 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_105_2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_4_247 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_122_602 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_107_698 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_106_164 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_121_134 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_96_34 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_453 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
Xhold50 hold50/I hold50/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
XFILLER_76_744 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_486 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_48_424 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xhold83 hold83/I hold83/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
Xhold61 hold61/I hold61/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
Xhold72 hold72/I hold72/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
XFILLER_102_392 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xhold94 hold94/I hold94/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
XFILLER_29_682 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_91_769 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_63_449 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_16_310 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_16_321 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_71_460 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_177_808 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_71_482 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_71_471 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_43_195 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XPHY_360 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_176_318 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_31_357 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_129_223 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_129_212 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_61_70 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_8_531 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_177_70 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4360_ _7902_/Q _4360_/A2 _7435_/Q _6623_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_4291_ _7973_/Q _4291_/A2 _4291_/B _4292_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi21_2
XFILLER_140_443 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_98_335 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_140_454 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6030_ hold64/Z _6038_/A2 _6030_/B _7655_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_101_808 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_98_379 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_100_318 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xclkbuf_0__1040_ _4036_/ZN clkbuf_0__1040_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XTAP_368 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_379 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_20_2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_39_424 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_66_254 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_67_799 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_66_265 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_82_747 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_81_224 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6932_ _7914_/Q _7913_/Q _6937_/A1 _6950_/A1 _7195_/C1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor4_4
XPHY_19 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_35_641 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_62_460 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6863_ _7504_/Q _6885_/A2 _6893_/B1 _7389_/Q _6864_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_5814_ _6539_/A1 _5816_/A2 _5814_/B hold777/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_167_318 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6794_ _7705_/Q _6889_/A2 _6894_/C1 _7835_/Q _6800_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_5745_ _5579_/B _5804_/A2 _5766_/A2 _5744_/Z _5747_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor4_1
XFILLER_50_688 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5676_ _5747_/A1 _5676_/A2 _5748_/A1 _5676_/B2 _5719_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai22_1
X_4627_ _7451_/Q _3830_/Z _4627_/B hold569/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_163_524 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7415_ _7415_/D _7306_/Z _4398_/I1 _7415_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_135_215 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xhold520 _7464_/Q hold520/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
XFILLER_151_708 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_135_248 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7346_ _7346_/D _7301_/Z _4415_/A2 _7346_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
Xhold531 hold531/I _7442_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
XFILLER_144_760 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_104_602 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xhold542 _7680_/Q hold542/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
Xhold553 _7656_/Q hold553/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
XFILLER_2_729 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4558_ _4454_/Z _4558_/A2 _4558_/B _7386_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_7277_ _7277_/A1 _7280_/A2 _7277_/B _7277_/C _7278_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi211_1
Xhold564 _7450_/Q hold564/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
Xhold575 _7710_/Q hold575/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
XFILLER_143_292 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_131_432 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_106_11 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
Xhold586 _7856_/Q hold586/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
X_4489_ hold841/Z _4504_/A2 hold842/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
Xhold597 _7523_/Q hold597/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
X_6228_ hold47/Z hold6/Z _6228_/B _7748_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_106_33 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_103_167 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_89_357 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6159_ hold488/Z _6174_/A2 _6160_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_880 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_106_88 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_66_59 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_66_37 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_891 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_57_221 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_122_21 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_85_574 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_72_246 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_122_76 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_82_69 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_81_780 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_13_302 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_25_173 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_26_685 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_158_318 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_13_357 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_40_176 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_182_811 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_181_354 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_31_73 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_147_73 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_5_567 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_134_281 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_134_270 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_110_605 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xinput140 wb_dat_i[20] _7259_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyb_1
Xinput162 wb_sel_i[1] _7281_/C2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyb_1
Xinput151 wb_dat_i[30] _7270_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XFILLER_49_777 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_48_287 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_64_747 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_17_641 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_44_460 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3860_ hold72/Z hold82/Z _6367_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_4
XFILLER_16_195 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_177_638 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_176_126 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3791_ _7336_/Q _4383_/A1 _4323_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_5530_ _5548_/A2 _5540_/B2 _5530_/B _5803_/A4 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XPHY_190 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
X_5461_ _5461_/A1 _5461_/A2 _5460_/Z _5461_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__and3_1
XFILLER_117_215 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_172_354 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_172_321 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4412_ _7441_/Q input93/Z _7585_/Q _4412_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_117_248 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_68_2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7200_ _7394_/Q _7200_/A2 _7200_/B1 _7388_/Q _7206_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_5392_ _5392_/A1 _5392_/A2 _5376_/B _5405_/B _5392_/B2 _5581_/C VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai32_1
X_4343_ _7520_/Q _4438_/A2 _7515_/Q _4344_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_125_281 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_113_421 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_7131_ _7433_/Q _7936_/Q _7132_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_7062_ _7858_/Q _6938_/I _7188_/A2 _7379_/Q _7063_/A4 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_4274_ _4274_/A1 _4274_/A2 _4274_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_101_649 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_101_638 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_100_104 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_98_187 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6013_ hold64/Z _6021_/A2 _6013_/B _7647_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_67_541 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_55_714 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7964_ _7964_/D _7317_/Z _4398_/I1 _7964_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XTAP_1309 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_6915_ _6937_/A1 _6953_/A1 _6599_/Z _7197_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor3_4
XFILLER_42_419 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_23_611 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_23_633 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_7895_ _7895_/D _7900_/RN _7900_/CLK _7895_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_168_605 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_167_104 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6846_ _7755_/Q _6644_/Z _6885_/B1 _7715_/Q _6847_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_11_806 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6777_ _6777_/A1 _6777_/A2 _6777_/A3 _6778_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor3_1
XFILLER_22_176 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_23_688 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_50_463 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_5728_ _5287_/C _5316_/B _5762_/A4 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_3989_ _3989_/A1 _3989_/A2 _3989_/A3 _3989_/A4 _3990_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand4_1
XFILLER_182_107 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_176_671 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5659_ _5674_/A1 _5674_/A2 _5657_/Z _5674_/A3 _5675_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand4_1
XFILLER_163_354 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_2_515 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7329_ _7901_/RN _4334_/Z _7329_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__and2_1
Xhold350 _7737_/Q hold350/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
Xhold361 hold361/I _4504_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
Xhold383 hold383/I _7428_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
Xhold372 _7795_/Q hold372/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
XFILLER_89_154 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
Xhold394 hold394/I _4895_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
XFILLER_93_24 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_46_703 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_172_2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_133_86 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_46_747 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1843 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1832 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1821 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1810 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_60_238 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_26_460 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1876 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1865 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1854 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1898 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1887 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_13_165 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_41_496 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_6_810 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_154_321 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_115_708 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_142_505 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_108_760 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_154_398 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_123_774 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_107_292 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_1_570 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_3_33 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_3_99 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_49_574 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_64_566 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4961_ _5022_/B _4944_/Z _4963_/A4 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_45_780 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3912_ _7691_/Q _6090_/A1 hold90/I _7723_/Q _3916_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_7680_ _7680_/D _7923_/RN _7737_/CLK _7680_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
X_4892_ _4454_/Z _4892_/A2 _4892_/B _7536_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_6700_ _7717_/Q _6881_/A2 _6882_/B1 _7653_/Q _6702_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_3843_ _3801_/Z _3864_/A2 _3843_/A3 _3864_/A4 _4075_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand4_4
XFILLER_32_463 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6631_ _7909_/Q _7908_/Q _6662_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_4
XFILLER_149_159 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_158_660 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3774_ _7345_/Q _3774_/A2 _3763_/B _3774_/B _7965_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai31_1
XFILLER_118_524 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_6562_ _6562_/A1 _6561_/Z _6564_/B _6563_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_173_641 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6493_ hold458/Z _6502_/A2 hold459/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_5513_ _5179_/B _5793_/A2 _5555_/B _5514_/A4 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_172_140 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_145_376 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_145_354 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5444_ _5627_/A2 _5444_/A2 _5613_/A2 _5444_/A4 _5445_/A4 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand4_1
XFILLER_154_19 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5375_ _5015_/B _5197_/Z _5375_/A3 _5375_/A4 _5708_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor4_4
X_7114_ _7900_/Q _7197_/A2 _7196_/A2 _7892_/Q _7196_/B1 _7642_/Q _7116_/A3 VDD VSS
+ gf180mcu_fd_sc_mcu7t5v0__aoi222_1
X_4326_ _7411_/Q _3738_/Z _4327_/S VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_141_560 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_99_496 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7045_ _7761_/Q _7202_/C2 _7205_/A2 _7735_/Q _7048_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_75_809 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4257_ _7504_/Q _4831_/A1 _5852_/A1 _4215_/Z _4260_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_86_179 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4188_ _7863_/Q _6469_/A1 _4554_/A1 _7386_/Q _7356_/Q _4488_/A1 _4203_/A2 VDD VSS
+ gf180mcu_fd_sc_mcu7t5v0__aoi222_2
XFILLER_28_747 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_103_45 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_103_56 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_103_89 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_7947_ _7947_/D _7949_/CLK _7947_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_70_536 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1117 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1128 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1106 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_27_279 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_43_739 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_70_547 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1139 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_7878_ _7878_/D _7900_/RN _7878_/CLK _7878_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffsnq_1
X_6829_ _7133_/S _6829_/A2 _6829_/B _7927_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_23_474 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_51_783 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_10_124 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_149_682 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_7_618 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_164_630 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_136_321 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_10_179 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_163_173 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_88_46 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_151_357 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_2_334 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xhold180 hold180/I _5996_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
Xhold191 hold191/I _7659_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
XFILLER_105_774 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_2_389 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_120_733 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_92_127 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_92_116 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_34_717 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_46_566 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2352 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2341 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2330 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2396 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2385 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2374 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2363 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1651 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1640 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1684 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1673 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1662 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_14_463 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_159_457 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1695 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_41_282 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_155_641 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_155_685 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_127_354 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_69_603 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_170_688 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5160_ _5538_/A1 _5390_/A2 _5162_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_5091_ _5058_/Z _5456_/A2 _5114_/A3 _5579_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__and3_2
XFILLER_110_210 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4111_ hold27/Z hold149/Z _5881_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_57_809 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4042_ _7793_/Q _6316_/A1 _4067_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_68_179 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_7801_ _7801_/D _7901_/RN _7833_/CLK _7801_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
X_5993_ hold596/Z _6004_/A2 _5994_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_4944_ _5338_/A1 _4900_/Z _4944_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__xor2_2
X_7732_ _7732_/D _7938_/RN _7791_/CLK _7732_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffsnq_1
XFILLER_33_783 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_178_766 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_177_232 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7663_ _7663_/D _7853_/RN _7726_/CLK hold79/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_20_433 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4875_ hold47/Z _4877_/A2 _4875_/B hold606/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_7594_ _7594_/D _7900_/RN _7897_/CLK _8004_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
X_3826_ hold76/Z hold38/Z _5954_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_4
X_6614_ _6953_/A2 _6950_/A2 _6955_/A4 _7193_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor3_4
X_3757_ _3765_/A1 _3765_/A2 _3762_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_118_321 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_6545_ _6545_/A1 _6553_/A2 _6545_/B hold178/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_173_471 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_173_482 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_161_611 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_133_302 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3688_ _7793_/Q _3688_/ZN VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_118_398 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6476_ hold98/Z _6485_/A2 hold99/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
Xoutput230 _8003_/Z mgmt_gpio_out[29] VDD VSS gf180mcu_fd_sc_mcu7t5v0__buf_4
XFILLER_133_357 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5427_ _5685_/B _5247_/B _5540_/C _5686_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi21_1
Xoutput252 _4422_/ZN pad_flash_io0_ie VDD VSS gf180mcu_fd_sc_mcu7t5v0__buf_4
Xoutput241 _7985_/Z mgmt_gpio_out[4] VDD VSS gf180mcu_fd_sc_mcu7t5v0__buf_4
XFILLER_160_176 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5358_ _5741_/A1 _5602_/A1 _5741_/A3 _5636_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor3_2
XFILLER_114_560 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
Xoutput274 _7359_/Q pll_trim[12] VDD VSS gf180mcu_fd_sc_mcu7t5v0__buf_4
Xoutput263 _7559_/Q pll_div[1] VDD VSS gf180mcu_fd_sc_mcu7t5v0__buf_4
Xoutput285 _7353_/Q pll_trim[22] VDD VSS gf180mcu_fd_sc_mcu7t5v0__buf_4
X_4309_ _4308_/Z _7340_/Q _4309_/S _7340_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_102_744 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_87_455 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xoutput296 _7356_/Q pll_trim[9] VDD VSS gf180mcu_fd_sc_mcu7t5v0__buf_4
X_5289_ _3723_/I _5579_/B _5721_/C _5680_/C _5293_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XFILLER_102_788 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_7028_ _7433_/Q _7932_/Q _7028_/B _7030_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_74_105 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_87_499 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_114_88 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_114_77 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_74_37 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_43_514 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_130_54 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_169_733 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_168_210 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_90_25 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_23_282 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_135_2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_139_63 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_137_641 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_128_129 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_11_499 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_152_600 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_139_85 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_109_354 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_109_343 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_152_666 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_155_73 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_152_688 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_151_176 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_709 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_93_425 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_78_499 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_19_544 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_80_108 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_74_672 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_62_812 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2171 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2160 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_34_547 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2193 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2182 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
Xnet299_2 net299_2/I _4416_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_15_761 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_159_232 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1492 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1481 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1470 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_14_271 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_15_783 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_30_731 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_174_202 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4660_ hold618/Z _3879_/Z _4660_/B _4661_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_147_438 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6330_ _4481_/I _6332_/A2 _6330_/B _7796_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_4591_ _6539_/A1 _4593_/A2 _4591_/B _7399_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_143_611 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_115_313 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xhold905 hold905/I _5816_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
Xhold927 _7348_/Q hold927/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
Xhold916 _7733_/Q hold916/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
XFILLER_50_2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xhold938 _7953_/Q _3670_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
X_6261_ hold378/Z _6264_/A2 hold379/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_115_357 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_89_709 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xhold949 _7552_/Q hold949/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
XFILLER_170_463 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5212_ _4906_/Z _5373_/A3 _5373_/A4 _5212_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__and3_1
XFILLER_142_176 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_142_154 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_8000_ _8000_/I _8000_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_6192_ _6192_/A1 _7285_/A2 _6208_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_4
X_5143_ _5645_/A1 _5545_/A2 _5768_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_142_198 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_97_753 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_97_775 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_28_19 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5074_ _5600_/A1 _5797_/B _5783_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_4
XFILLER_111_596 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_84_436 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_84_425 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_69_499 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_56_105 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_56_138 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4025_ _4025_/A1 _4025_/A2 _4025_/A3 _4025_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__or3_1
XFILLER_72_609 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_80_631 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5976_ hold687/Z _5987_/A2 _5977_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_13_709 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4927_ _5211_/A3 _4920_/Z _5011_/B _4951_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi21_2
X_7715_ _7715_/D _7853_/RN _7812_/CLK _7715_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_33_580 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_7646_ _7646_/D _7961_/RN _7650_/CLK _7646_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffsnq_1
XFILLER_20_241 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4858_ _4858_/A1 _7285_/A2 _4862_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_166_747 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_165_224 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3809_ hold49/Z hold80/Z _3811_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_20_263 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_21_775 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_119_641 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_109_11 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7577_ _7577_/D _7961_/RN _7624_/CLK _7577_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
X_4789_ _7480_/Q _4795_/S _4790_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_181_739 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_146_471 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_146_460 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_119_685 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_109_44 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_109_33 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6528_ _6545_/A1 _6536_/A2 _6528_/B hold172/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_161_441 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_118_195 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6459_ hold160/Z _6468_/A2 hold161/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
Xclkbuf_leaf_7_csclk clkbuf_leaf_9_csclk/I _7866_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_161_496 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_102_563 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_102_552 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_85_58 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_75_425 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_28_330 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_141_64 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_62_108 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_44_812 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_55_160 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_56_672 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_141_97 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_70_130 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_169_552 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_34_51 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_43_399 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_156_202 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_12_742 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_7_212 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_172_717 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_109_140 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_125_611 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_152_463 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_124_176 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_506 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_59_70 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_539 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_528 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_517 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_78_241 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_66_425 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_38_105 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_54_609 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_81_439 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_81_428 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_35_812 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_179_305 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_34_311 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_61_141 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5830_ _6539_/A1 _5840_/A2 _5830_/B _7563_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_5761_ _5686_/Z _5761_/A2 _5758_/Z _5760_/Z _5786_/B1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand4_1
XFILLER_98_2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4712_ _3819_/Z _4481_/I _4713_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_7500_ _7500_/D _7949_/CLK _7500_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_148_747 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_147_235 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5692_ _5692_/A1 _5692_/A2 _5692_/B _5694_/A4 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_7431_ _7431_/D _7923_/RN _7597_/CLK _7987_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_147_246 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4643_ _7455_/Q _3830_/Z _4643_/B _4644_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_128_460 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xhold702 hold702/I _6121_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
X_7362_ _7362_/D input75/Z _7875_/CLK _7362_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffsnq_1
X_4574_ _4574_/A1 _6537_/A2 _4578_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_7293_ _7901_/RN _4334_/Z _7293_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_155_290 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_115_121 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
Xhold724 _7641_/Q hold724/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
X_6313_ hold233/Z _6315_/A2 _6313_/B hold308/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
Xhold713 hold713/I _6087_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
Xhold746 hold746/I _4500_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
Xhold735 _7531_/Q hold735/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
XFILLER_171_783 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_171_761 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_115_176 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xhold757 _7395_/Q hold757/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
Xhold779 _7466_/Q hold779/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
Xhold768 _7535_/Q hold768/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
X_6244_ hold748/Z _6247_/A2 _6245_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_170_282 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_143_496 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_131_636 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_131_647 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_6175_ hold28/Z _7285_/A2 _6191_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_4
XFILLER_85_712 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_57_403 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5126_ _5390_/A2 _5122_/Z _5479_/A2 _5669_/A1 _5651_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_130_179 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_57_414 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_57_436 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5057_ _5303_/A3 _5421_/A1 _5319_/C VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_4
XFILLER_84_244 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_55_17 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_57_458 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4008_ _7624_/Q _5954_/A1 _4020_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_25_300 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_26_812 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_38_672 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_44_108 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_25_366 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_53_664 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_53_653 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5959_ hold582/Z _5970_/A2 _5960_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_139_714 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_40_347 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_21_550 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7629_ _7629_/D _7877_/RN _7752_/CLK _7629_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffsnq_1
XFILLER_147_780 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_181_558 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_107_655 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_134_463 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_136_75 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_106_176 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_96_13 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_96_46 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
Xhold40 hold40/I hold40/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
Xhold62 hold62/I hold62/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
Xhold51 hold51/I hold51/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
Xhold73 hold73/I hold73/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
XFILLER_152_52 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_75_233 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_29_73 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_152_96 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
Xhold84 hold84/I hold84/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
Xhold95 hold95/I hold95/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
XFILLER_63_428 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_17_812 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_90_247 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_29_694 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_16_366 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_43_141 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_71_494 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_16_388 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_43_185 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_361 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_350 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_61_82 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_172_514 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_145_728 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_144_205 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_8_587 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_6_33 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_125_430 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_153_783 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_125_452 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_4290_ _7973_/Q _4291_/A2 _4382_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_152_271 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_125_496 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_98_325 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_140_488 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_112_179 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_67_712 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_369 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_94_531 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_13_2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_7980_ _7980_/D _7333_/Z _4398_/I1 _7980_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_26_108 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_6931_ _6937_/A1 _6941_/A1 _7196_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_4
XFILLER_34_141 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6862_ _7405_/Q _6883_/A2 _6883_/B1 _7397_/Q _6864_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_5813_ hold775/Z _5816_/A2 hold776/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_6793_ _7641_/Q _6890_/A2 _6665_/Z _7745_/Q _6793_/C _6800_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi221_1
X_5744_ _5499_/Z _5542_/Z _5744_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__or2_1
XFILLER_148_544 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_136_717 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_5675_ _5675_/A1 _5671_/Z _5676_/B2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_1
Xclkbuf_leaf_72_csclk clkbuf_3_3__f_csclk/Z _7741_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
X_4626_ _3830_/Z _4454_/Z hold568/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_7414_ _7414_/D _7305_/Z _4415_/A2 _7414_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_4
XFILLER_135_227 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_129_780 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7345_ _7345_/D _7300_/Z _4398_/I1 _7345_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_2
XFILLER_135_238 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
Xhold510 _7674_/Q hold510/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
Xhold521 hold521/I hold521/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
XFILLER_116_463 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xhold543 hold543/I _6083_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
Xhold554 _7736_/Q hold554/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
Xhold532 _7565_/Q hold532/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
X_4557_ hold869/Z _4558_/A2 _4558_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_7276_ _7276_/A1 _7276_/A2 _7277_/C VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
Xhold565 hold565/I hold565/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
Xhold576 hold576/I _6147_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
XFILLER_104_625 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_89_347 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
Xclkbuf_leaf_87_csclk _7528_/CLK _7627_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
X_4488_ _4488_/A1 _6537_/A2 _4504_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_4
Xhold587 _7468_/Q hold587/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
X_6227_ hold486/Z hold6/Z _6228_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
Xhold598 hold598/I _4860_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
XFILLER_131_499 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_6158_ hold90/Z _7285_/A2 _6174_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_4
XFILLER_106_78 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_870 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_58_734 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5109_ _5669_/A1 _5672_/A2 _5673_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_85_531 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_881 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_892 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
Xclkbuf_leaf_10_csclk clkbuf_leaf_9_csclk/I _7830_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
X_6089_ _6553_/A1 _6089_/A2 _6089_/B hold186/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_73_737 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_45_428 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xclkbuf_leaf_25_csclk _7422_/CLK _7877_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_122_88 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_122_66 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_82_37 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_14_804 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_25_141 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_25_163 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_53_472 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_40_133 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_41_667 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_139_555 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_127_706 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_40_188 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_154_514 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_154_558 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_147_85 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_135_783 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_107_474 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_107_463 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_122_400 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_107_496 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_107_485 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_163_73 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_49_712 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xinput152 wb_dat_i[31] _7275_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyb_1
Xinput130 wb_dat_i[11] _7255_/B1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyb_1
Xinput141 wb_dat_i[21] _7265_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyb_1
Xinput163 wb_sel_i[2] _7281_/B1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XFILLER_102_190 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_76_531 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_76_542 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_76_520 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_91_567 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_63_269 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_72_770 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_176_105 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_20_807 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3790_ hold74/Z _3789_/Z _3810_/S hold75/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_4
XFILLER_31_144 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_191 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_180 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_173_812 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_172_300 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_145_503 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5460_ _5460_/A1 _5460_/A2 _5657_/A3 _5460_/A4 _5460_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__and4_1
XFILLER_172_333 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4411_ _7442_/Q _4411_/I1 _7583_/Q _4411_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_133_709 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_132_208 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5391_ _5741_/A1 _4993_/B _5797_/A1 _5391_/B _5735_/C VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai31_1
X_4342_ _4342_/I _7519_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_7130_ _7130_/A1 _7130_/A2 _7130_/A3 _6949_/I _7610_/Q _7132_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai32_1
X_7061_ _7648_/Q _7195_/A2 _7195_/B1 _7624_/Q _7195_/C1 _7874_/Q _7063_/A3 VDD VSS
+ gf180mcu_fd_sc_mcu7t5v0__aoi222_1
X_4273_ _7563_/Q hold150/I _4574_/A1 _7393_/Q _4274_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_113_499 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6012_ hold78/Z _6021_/A2 _6013_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
.ends

