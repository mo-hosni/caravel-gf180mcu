magic
tech gf180mcuC
magscale 1 10
timestamp 1668683681
<< metal1 >>
rect 224 10218 16688 10252
rect 224 10166 2152 10218
rect 2204 10166 2256 10218
rect 2308 10166 2360 10218
rect 2412 10166 6268 10218
rect 6320 10166 6372 10218
rect 6424 10166 6476 10218
rect 6528 10166 10384 10218
rect 10436 10166 10488 10218
rect 10540 10166 10592 10218
rect 10644 10166 14500 10218
rect 14552 10166 14604 10218
rect 14656 10166 14708 10218
rect 14760 10166 16688 10218
rect 224 10132 16688 10166
rect 15486 9938 15538 9950
rect 1474 9886 1486 9938
rect 1538 9886 1550 9938
rect 13906 9886 13918 9938
rect 13970 9886 13982 9938
rect 15486 9874 15538 9886
rect 3378 9774 3390 9826
rect 3442 9774 3454 9826
rect 14914 9774 14926 9826
rect 14978 9774 14990 9826
rect 4622 9602 4674 9614
rect 4622 9538 4674 9550
rect 5070 9602 5122 9614
rect 5070 9538 5122 9550
rect 224 9434 16848 9468
rect 224 9382 4210 9434
rect 4262 9382 4314 9434
rect 4366 9382 4418 9434
rect 4470 9382 8326 9434
rect 8378 9382 8430 9434
rect 8482 9382 8534 9434
rect 8586 9382 12442 9434
rect 12494 9382 12546 9434
rect 12598 9382 12650 9434
rect 12702 9382 16558 9434
rect 16610 9382 16662 9434
rect 16714 9382 16766 9434
rect 16818 9382 16848 9434
rect 224 9348 16848 9382
rect 15486 9042 15538 9054
rect 4386 8990 4398 9042
rect 4450 8990 4462 9042
rect 5282 8990 5294 9042
rect 5346 8990 5358 9042
rect 11666 8990 11678 9042
rect 11730 8990 11742 9042
rect 14466 8990 14478 9042
rect 14530 8990 14542 9042
rect 15486 8978 15538 8990
rect 2818 8878 2830 8930
rect 2882 8878 2894 8930
rect 7634 8878 7646 8930
rect 7698 8878 7710 8930
rect 10770 8878 10782 8930
rect 10834 8878 10846 8930
rect 13906 8878 13918 8930
rect 13970 8878 13982 8930
rect 224 8650 16688 8684
rect 224 8598 2152 8650
rect 2204 8598 2256 8650
rect 2308 8598 2360 8650
rect 2412 8598 6268 8650
rect 6320 8598 6372 8650
rect 6424 8598 6476 8650
rect 6528 8598 10384 8650
rect 10436 8598 10488 8650
rect 10540 8598 10592 8650
rect 10644 8598 14500 8650
rect 14552 8598 14604 8650
rect 14656 8598 14708 8650
rect 14760 8598 16688 8650
rect 224 8564 16688 8598
rect 5070 8370 5122 8382
rect 11902 8370 11954 8382
rect 1922 8318 1934 8370
rect 1986 8318 1998 8370
rect 7746 8318 7758 8370
rect 7810 8318 7822 8370
rect 13458 8318 13470 8370
rect 13522 8318 13534 8370
rect 5070 8306 5122 8318
rect 11902 8306 11954 8318
rect 15598 8258 15650 8270
rect 3490 8206 3502 8258
rect 3554 8206 3566 8258
rect 8866 8206 8878 8258
rect 8930 8206 8942 8258
rect 14578 8206 14590 8258
rect 14642 8206 14654 8258
rect 15598 8194 15650 8206
rect 4510 8034 4562 8046
rect 4510 7970 4562 7982
rect 9886 8034 9938 8046
rect 9886 7970 9938 7982
rect 224 7866 16848 7900
rect 224 7814 4210 7866
rect 4262 7814 4314 7866
rect 4366 7814 4418 7866
rect 4470 7814 8326 7866
rect 8378 7814 8430 7866
rect 8482 7814 8534 7866
rect 8586 7814 12442 7866
rect 12494 7814 12546 7866
rect 12598 7814 12650 7866
rect 12702 7814 16558 7866
rect 16610 7814 16662 7866
rect 16714 7814 16766 7866
rect 16818 7814 16848 7866
rect 224 7780 16848 7814
rect 14142 7698 14194 7710
rect 14142 7634 14194 7646
rect 3714 7422 3726 7474
rect 3778 7422 3790 7474
rect 6290 7422 6302 7474
rect 6354 7422 6366 7474
rect 13122 7422 13134 7474
rect 13186 7422 13198 7474
rect 7310 7362 7362 7374
rect 2594 7310 2606 7362
rect 2658 7310 2670 7362
rect 5170 7310 5182 7362
rect 5234 7310 5246 7362
rect 12226 7310 12238 7362
rect 12290 7310 12302 7362
rect 7310 7298 7362 7310
rect 224 7082 16688 7116
rect 224 7030 2152 7082
rect 2204 7030 2256 7082
rect 2308 7030 2360 7082
rect 2412 7030 6268 7082
rect 6320 7030 6372 7082
rect 6424 7030 6476 7082
rect 6528 7030 10384 7082
rect 10436 7030 10488 7082
rect 10540 7030 10592 7082
rect 10644 7030 14500 7082
rect 14552 7030 14604 7082
rect 14656 7030 14708 7082
rect 14760 7030 16688 7082
rect 224 6996 16688 7030
rect 2482 6750 2494 6802
rect 2546 6750 2558 6802
rect 8194 6750 8206 6802
rect 8258 6750 8270 6802
rect 13122 6750 13134 6802
rect 13186 6750 13198 6802
rect 5406 6690 5458 6702
rect 11790 6690 11842 6702
rect 15598 6690 15650 6702
rect 3378 6638 3390 6690
rect 3442 6638 3454 6690
rect 9314 6638 9326 6690
rect 9378 6638 9390 6690
rect 14578 6638 14590 6690
rect 14642 6638 14654 6690
rect 5406 6626 5458 6638
rect 11790 6626 11842 6638
rect 15598 6626 15650 6638
rect 10334 6578 10386 6590
rect 10334 6514 10386 6526
rect 4510 6466 4562 6478
rect 4510 6402 4562 6414
rect 4958 6466 5010 6478
rect 4958 6402 5010 6414
rect 224 6298 16848 6332
rect 224 6246 4210 6298
rect 4262 6246 4314 6298
rect 4366 6246 4418 6298
rect 4470 6246 8326 6298
rect 8378 6246 8430 6298
rect 8482 6246 8534 6298
rect 8586 6246 12442 6298
rect 12494 6246 12546 6298
rect 12598 6246 12650 6298
rect 12702 6246 16558 6298
rect 16610 6246 16662 6298
rect 16714 6246 16766 6298
rect 16818 6246 16848 6298
rect 224 6212 16848 6246
rect 4162 5854 4174 5906
rect 4226 5854 4238 5906
rect 7522 5854 7534 5906
rect 7586 5854 7598 5906
rect 10994 5854 11006 5906
rect 11058 5854 11070 5906
rect 12114 5854 12126 5906
rect 12178 5854 12190 5906
rect 3042 5742 3054 5794
rect 3106 5742 3118 5794
rect 6626 5742 6638 5794
rect 6690 5742 6702 5794
rect 9986 5742 9998 5794
rect 10050 5742 10062 5794
rect 13682 5742 13694 5794
rect 13746 5742 13758 5794
rect 224 5514 16688 5548
rect 224 5462 2152 5514
rect 2204 5462 2256 5514
rect 2308 5462 2360 5514
rect 2412 5462 6268 5514
rect 6320 5462 6372 5514
rect 6424 5462 6476 5514
rect 6528 5462 10384 5514
rect 10436 5462 10488 5514
rect 10540 5462 10592 5514
rect 10644 5462 14500 5514
rect 14552 5462 14604 5514
rect 14656 5462 14708 5514
rect 14760 5462 16688 5514
rect 224 5428 16688 5462
rect 11790 5234 11842 5246
rect 15598 5234 15650 5246
rect 2706 5182 2718 5234
rect 2770 5182 2782 5234
rect 5954 5182 5966 5234
rect 6018 5182 6030 5234
rect 9538 5182 9550 5234
rect 9602 5182 9614 5234
rect 14018 5182 14030 5234
rect 14082 5182 14094 5234
rect 11790 5170 11842 5182
rect 15598 5170 15650 5182
rect 4510 5122 4562 5134
rect 3826 5070 3838 5122
rect 3890 5070 3902 5122
rect 7186 5070 7198 5122
rect 7250 5070 7262 5122
rect 10770 5070 10782 5122
rect 10834 5070 10846 5122
rect 15026 5070 15038 5122
rect 15090 5070 15102 5122
rect 4510 5058 4562 5070
rect 224 4730 16848 4764
rect 224 4678 4210 4730
rect 4262 4678 4314 4730
rect 4366 4678 4418 4730
rect 4470 4678 8326 4730
rect 8378 4678 8430 4730
rect 8482 4678 8534 4730
rect 8586 4678 12442 4730
rect 12494 4678 12546 4730
rect 12598 4678 12650 4730
rect 12702 4678 16558 4730
rect 16610 4678 16662 4730
rect 16714 4678 16766 4730
rect 16818 4678 16848 4730
rect 224 4644 16848 4678
rect 7870 4562 7922 4574
rect 7870 4498 7922 4510
rect 8990 4562 9042 4574
rect 8990 4498 9042 4510
rect 1474 4398 1486 4450
rect 1538 4398 1550 4450
rect 6862 4338 6914 4350
rect 13694 4338 13746 4350
rect 3266 4286 3278 4338
rect 3330 4286 3342 4338
rect 5842 4286 5854 4338
rect 5906 4286 5918 4338
rect 12674 4286 12686 4338
rect 12738 4286 12750 4338
rect 6862 4274 6914 4286
rect 13694 4274 13746 4286
rect 8542 4226 8594 4238
rect 14142 4226 14194 4238
rect 4722 4174 4734 4226
rect 4786 4174 4798 4226
rect 11890 4174 11902 4226
rect 11954 4174 11966 4226
rect 8542 4162 8594 4174
rect 14142 4162 14194 4174
rect 224 3946 16688 3980
rect 224 3894 2152 3946
rect 2204 3894 2256 3946
rect 2308 3894 2360 3946
rect 2412 3894 6268 3946
rect 6320 3894 6372 3946
rect 6424 3894 6476 3946
rect 6528 3894 10384 3946
rect 10436 3894 10488 3946
rect 10540 3894 10592 3946
rect 10644 3894 14500 3946
rect 14552 3894 14604 3946
rect 14656 3894 14708 3946
rect 14760 3894 16688 3946
rect 224 3860 16688 3894
rect 15362 3726 15374 3778
rect 15426 3775 15438 3778
rect 16034 3775 16046 3778
rect 15426 3729 16046 3775
rect 15426 3726 15438 3729
rect 16034 3726 16046 3729
rect 16098 3726 16110 3778
rect 16046 3666 16098 3678
rect 2370 3614 2382 3666
rect 2434 3614 2446 3666
rect 6514 3614 6526 3666
rect 6578 3614 6590 3666
rect 9090 3614 9102 3666
rect 9154 3614 9166 3666
rect 10770 3614 10782 3666
rect 10834 3663 10846 3666
rect 11218 3663 11230 3666
rect 10834 3617 11230 3663
rect 10834 3614 10846 3617
rect 11218 3614 11230 3617
rect 11282 3614 11294 3666
rect 13570 3614 13582 3666
rect 13634 3614 13646 3666
rect 16046 3602 16098 3614
rect 11342 3554 11394 3566
rect 1250 3502 1262 3554
rect 1314 3502 1326 3554
rect 7634 3502 7646 3554
rect 7698 3502 7710 3554
rect 10210 3502 10222 3554
rect 10274 3502 10286 3554
rect 11342 3490 11394 3502
rect 11790 3554 11842 3566
rect 15598 3554 15650 3566
rect 14578 3502 14590 3554
rect 14642 3502 14654 3554
rect 11790 3490 11842 3502
rect 15598 3490 15650 3502
rect 702 3442 754 3454
rect 702 3378 754 3390
rect 4510 3442 4562 3454
rect 4510 3378 4562 3390
rect 224 3162 16848 3196
rect 224 3110 4210 3162
rect 4262 3110 4314 3162
rect 4366 3110 4418 3162
rect 4470 3110 8326 3162
rect 8378 3110 8430 3162
rect 8482 3110 8534 3162
rect 8586 3110 12442 3162
rect 12494 3110 12546 3162
rect 12598 3110 12650 3162
rect 12702 3110 16558 3162
rect 16610 3110 16662 3162
rect 16714 3110 16766 3162
rect 16818 3110 16848 3162
rect 224 3076 16848 3110
rect 1598 2994 1650 3006
rect 1598 2930 1650 2942
rect 6066 2830 6078 2882
rect 6130 2830 6142 2882
rect 8542 2770 8594 2782
rect 2146 2718 2158 2770
rect 2210 2718 2222 2770
rect 7298 2718 7310 2770
rect 7362 2718 7374 2770
rect 12002 2718 12014 2770
rect 12066 2718 12078 2770
rect 15474 2718 15486 2770
rect 15538 2718 15550 2770
rect 8542 2706 8594 2718
rect 4498 2606 4510 2658
rect 4562 2606 4574 2658
rect 10882 2606 10894 2658
rect 10946 2606 10958 2658
rect 14466 2606 14478 2658
rect 14530 2606 14542 2658
rect 224 2378 16688 2412
rect 224 2326 2152 2378
rect 2204 2326 2256 2378
rect 2308 2326 2360 2378
rect 2412 2326 6268 2378
rect 6320 2326 6372 2378
rect 6424 2326 6476 2378
rect 6528 2326 10384 2378
rect 10436 2326 10488 2378
rect 10540 2326 10592 2378
rect 10644 2326 14500 2378
rect 14552 2326 14604 2378
rect 14656 2326 14708 2378
rect 14760 2326 16688 2378
rect 224 2292 16688 2326
rect 15598 2098 15650 2110
rect 2482 2046 2494 2098
rect 2546 2046 2558 2098
rect 5506 2046 5518 2098
rect 5570 2046 5582 2098
rect 8754 2046 8766 2098
rect 8818 2046 8830 2098
rect 11106 2046 11118 2098
rect 11170 2095 11182 2098
rect 11442 2095 11454 2098
rect 11170 2049 11454 2095
rect 11170 2046 11182 2049
rect 11442 2046 11454 2049
rect 11506 2046 11518 2098
rect 13906 2046 13918 2098
rect 13970 2046 13982 2098
rect 15598 2034 15650 2046
rect 814 1986 866 1998
rect 11566 1986 11618 1998
rect 1250 1934 1262 1986
rect 1314 1934 1326 1986
rect 6738 1934 6750 1986
rect 6802 1934 6814 1986
rect 11106 1934 11118 1986
rect 11170 1934 11182 1986
rect 15026 1934 15038 1986
rect 15090 1934 15102 1986
rect 814 1922 866 1934
rect 11566 1922 11618 1934
rect 7758 1874 7810 1886
rect 7758 1810 7810 1822
rect 224 1594 16848 1628
rect 224 1542 4210 1594
rect 4262 1542 4314 1594
rect 4366 1542 4418 1594
rect 4470 1542 8326 1594
rect 8378 1542 8430 1594
rect 8482 1542 8534 1594
rect 8586 1542 12442 1594
rect 12494 1542 12546 1594
rect 12598 1542 12650 1594
rect 12702 1542 16558 1594
rect 16610 1542 16662 1594
rect 16714 1542 16766 1594
rect 16818 1542 16848 1594
rect 224 1508 16848 1542
<< via1 >>
rect 2152 10166 2204 10218
rect 2256 10166 2308 10218
rect 2360 10166 2412 10218
rect 6268 10166 6320 10218
rect 6372 10166 6424 10218
rect 6476 10166 6528 10218
rect 10384 10166 10436 10218
rect 10488 10166 10540 10218
rect 10592 10166 10644 10218
rect 14500 10166 14552 10218
rect 14604 10166 14656 10218
rect 14708 10166 14760 10218
rect 1486 9886 1538 9938
rect 13918 9886 13970 9938
rect 15486 9886 15538 9938
rect 3390 9774 3442 9826
rect 14926 9774 14978 9826
rect 4622 9550 4674 9602
rect 5070 9550 5122 9602
rect 4210 9382 4262 9434
rect 4314 9382 4366 9434
rect 4418 9382 4470 9434
rect 8326 9382 8378 9434
rect 8430 9382 8482 9434
rect 8534 9382 8586 9434
rect 12442 9382 12494 9434
rect 12546 9382 12598 9434
rect 12650 9382 12702 9434
rect 16558 9382 16610 9434
rect 16662 9382 16714 9434
rect 16766 9382 16818 9434
rect 4398 8990 4450 9042
rect 5294 8990 5346 9042
rect 11678 8990 11730 9042
rect 14478 8990 14530 9042
rect 15486 8990 15538 9042
rect 2830 8878 2882 8930
rect 7646 8878 7698 8930
rect 10782 8878 10834 8930
rect 13918 8878 13970 8930
rect 2152 8598 2204 8650
rect 2256 8598 2308 8650
rect 2360 8598 2412 8650
rect 6268 8598 6320 8650
rect 6372 8598 6424 8650
rect 6476 8598 6528 8650
rect 10384 8598 10436 8650
rect 10488 8598 10540 8650
rect 10592 8598 10644 8650
rect 14500 8598 14552 8650
rect 14604 8598 14656 8650
rect 14708 8598 14760 8650
rect 1934 8318 1986 8370
rect 5070 8318 5122 8370
rect 7758 8318 7810 8370
rect 11902 8318 11954 8370
rect 13470 8318 13522 8370
rect 3502 8206 3554 8258
rect 8878 8206 8930 8258
rect 14590 8206 14642 8258
rect 15598 8206 15650 8258
rect 4510 7982 4562 8034
rect 9886 7982 9938 8034
rect 4210 7814 4262 7866
rect 4314 7814 4366 7866
rect 4418 7814 4470 7866
rect 8326 7814 8378 7866
rect 8430 7814 8482 7866
rect 8534 7814 8586 7866
rect 12442 7814 12494 7866
rect 12546 7814 12598 7866
rect 12650 7814 12702 7866
rect 16558 7814 16610 7866
rect 16662 7814 16714 7866
rect 16766 7814 16818 7866
rect 14142 7646 14194 7698
rect 3726 7422 3778 7474
rect 6302 7422 6354 7474
rect 13134 7422 13186 7474
rect 2606 7310 2658 7362
rect 5182 7310 5234 7362
rect 7310 7310 7362 7362
rect 12238 7310 12290 7362
rect 2152 7030 2204 7082
rect 2256 7030 2308 7082
rect 2360 7030 2412 7082
rect 6268 7030 6320 7082
rect 6372 7030 6424 7082
rect 6476 7030 6528 7082
rect 10384 7030 10436 7082
rect 10488 7030 10540 7082
rect 10592 7030 10644 7082
rect 14500 7030 14552 7082
rect 14604 7030 14656 7082
rect 14708 7030 14760 7082
rect 2494 6750 2546 6802
rect 8206 6750 8258 6802
rect 13134 6750 13186 6802
rect 3390 6638 3442 6690
rect 5406 6638 5458 6690
rect 9326 6638 9378 6690
rect 11790 6638 11842 6690
rect 14590 6638 14642 6690
rect 15598 6638 15650 6690
rect 10334 6526 10386 6578
rect 4510 6414 4562 6466
rect 4958 6414 5010 6466
rect 4210 6246 4262 6298
rect 4314 6246 4366 6298
rect 4418 6246 4470 6298
rect 8326 6246 8378 6298
rect 8430 6246 8482 6298
rect 8534 6246 8586 6298
rect 12442 6246 12494 6298
rect 12546 6246 12598 6298
rect 12650 6246 12702 6298
rect 16558 6246 16610 6298
rect 16662 6246 16714 6298
rect 16766 6246 16818 6298
rect 4174 5854 4226 5906
rect 7534 5854 7586 5906
rect 11006 5854 11058 5906
rect 12126 5854 12178 5906
rect 3054 5742 3106 5794
rect 6638 5742 6690 5794
rect 9998 5742 10050 5794
rect 13694 5742 13746 5794
rect 2152 5462 2204 5514
rect 2256 5462 2308 5514
rect 2360 5462 2412 5514
rect 6268 5462 6320 5514
rect 6372 5462 6424 5514
rect 6476 5462 6528 5514
rect 10384 5462 10436 5514
rect 10488 5462 10540 5514
rect 10592 5462 10644 5514
rect 14500 5462 14552 5514
rect 14604 5462 14656 5514
rect 14708 5462 14760 5514
rect 2718 5182 2770 5234
rect 5966 5182 6018 5234
rect 9550 5182 9602 5234
rect 11790 5182 11842 5234
rect 14030 5182 14082 5234
rect 15598 5182 15650 5234
rect 3838 5070 3890 5122
rect 4510 5070 4562 5122
rect 7198 5070 7250 5122
rect 10782 5070 10834 5122
rect 15038 5070 15090 5122
rect 4210 4678 4262 4730
rect 4314 4678 4366 4730
rect 4418 4678 4470 4730
rect 8326 4678 8378 4730
rect 8430 4678 8482 4730
rect 8534 4678 8586 4730
rect 12442 4678 12494 4730
rect 12546 4678 12598 4730
rect 12650 4678 12702 4730
rect 16558 4678 16610 4730
rect 16662 4678 16714 4730
rect 16766 4678 16818 4730
rect 7870 4510 7922 4562
rect 8990 4510 9042 4562
rect 1486 4398 1538 4450
rect 3278 4286 3330 4338
rect 5854 4286 5906 4338
rect 6862 4286 6914 4338
rect 12686 4286 12738 4338
rect 13694 4286 13746 4338
rect 4734 4174 4786 4226
rect 8542 4174 8594 4226
rect 11902 4174 11954 4226
rect 14142 4174 14194 4226
rect 2152 3894 2204 3946
rect 2256 3894 2308 3946
rect 2360 3894 2412 3946
rect 6268 3894 6320 3946
rect 6372 3894 6424 3946
rect 6476 3894 6528 3946
rect 10384 3894 10436 3946
rect 10488 3894 10540 3946
rect 10592 3894 10644 3946
rect 14500 3894 14552 3946
rect 14604 3894 14656 3946
rect 14708 3894 14760 3946
rect 15374 3726 15426 3778
rect 16046 3726 16098 3778
rect 2382 3614 2434 3666
rect 6526 3614 6578 3666
rect 9102 3614 9154 3666
rect 10782 3614 10834 3666
rect 11230 3614 11282 3666
rect 13582 3614 13634 3666
rect 16046 3614 16098 3666
rect 1262 3502 1314 3554
rect 7646 3502 7698 3554
rect 10222 3502 10274 3554
rect 11342 3502 11394 3554
rect 11790 3502 11842 3554
rect 14590 3502 14642 3554
rect 15598 3502 15650 3554
rect 702 3390 754 3442
rect 4510 3390 4562 3442
rect 4210 3110 4262 3162
rect 4314 3110 4366 3162
rect 4418 3110 4470 3162
rect 8326 3110 8378 3162
rect 8430 3110 8482 3162
rect 8534 3110 8586 3162
rect 12442 3110 12494 3162
rect 12546 3110 12598 3162
rect 12650 3110 12702 3162
rect 16558 3110 16610 3162
rect 16662 3110 16714 3162
rect 16766 3110 16818 3162
rect 1598 2942 1650 2994
rect 6078 2830 6130 2882
rect 2158 2718 2210 2770
rect 7310 2718 7362 2770
rect 8542 2718 8594 2770
rect 12014 2718 12066 2770
rect 15486 2718 15538 2770
rect 4510 2606 4562 2658
rect 10894 2606 10946 2658
rect 14478 2606 14530 2658
rect 2152 2326 2204 2378
rect 2256 2326 2308 2378
rect 2360 2326 2412 2378
rect 6268 2326 6320 2378
rect 6372 2326 6424 2378
rect 6476 2326 6528 2378
rect 10384 2326 10436 2378
rect 10488 2326 10540 2378
rect 10592 2326 10644 2378
rect 14500 2326 14552 2378
rect 14604 2326 14656 2378
rect 14708 2326 14760 2378
rect 2494 2046 2546 2098
rect 5518 2046 5570 2098
rect 8766 2046 8818 2098
rect 11118 2046 11170 2098
rect 11454 2046 11506 2098
rect 13918 2046 13970 2098
rect 15598 2046 15650 2098
rect 814 1934 866 1986
rect 1262 1934 1314 1986
rect 6750 1934 6802 1986
rect 11118 1934 11170 1986
rect 11566 1934 11618 1986
rect 15038 1934 15090 1986
rect 7758 1822 7810 1874
rect 4210 1542 4262 1594
rect 4314 1542 4366 1594
rect 4418 1542 4470 1594
rect 8326 1542 8378 1594
rect 8430 1542 8482 1594
rect 8534 1542 8586 1594
rect 12442 1542 12494 1594
rect 12546 1542 12598 1594
rect 12650 1542 12702 1594
rect 16558 1542 16610 1594
rect 16662 1542 16714 1594
rect 16766 1542 16818 1594
<< metal2 >>
rect 560 11200 672 12000
rect 1008 11200 1120 12000
rect 1456 11200 1568 12000
rect 1904 11200 2016 12000
rect 2352 11200 2464 12000
rect 2800 11200 2912 12000
rect 3248 11200 3360 12000
rect 3696 11200 3808 12000
rect 4144 11200 4256 12000
rect 4592 11200 4704 12000
rect 5040 11200 5152 12000
rect 5488 11200 5600 12000
rect 5936 11200 6048 12000
rect 6384 11200 6496 12000
rect 6832 11200 6944 12000
rect 7280 11200 7392 12000
rect 7728 11200 7840 12000
rect 8176 11200 8288 12000
rect 8624 11200 8736 12000
rect 9072 11200 9184 12000
rect 9520 11200 9632 12000
rect 9968 11200 10080 12000
rect 10416 11200 10528 12000
rect 10864 11200 10976 12000
rect 11312 11200 11424 12000
rect 11760 11200 11872 12000
rect 12208 11200 12320 12000
rect 12656 11200 12768 12000
rect 13104 11200 13216 12000
rect 13552 11200 13664 12000
rect 14000 11200 14112 12000
rect 14448 11200 14560 12000
rect 14896 11200 15008 12000
rect 15344 11200 15456 12000
rect 15792 11200 15904 12000
rect 16240 11200 16352 12000
rect 588 3668 644 11200
rect 1036 5012 1092 11200
rect 1484 9938 1540 11200
rect 1484 9886 1486 9938
rect 1538 9886 1540 9938
rect 1484 9874 1540 9886
rect 1036 4946 1092 4956
rect 1596 9828 1652 9838
rect 1484 4452 1540 4462
rect 1484 4358 1540 4396
rect 1596 4004 1652 9772
rect 1932 8370 1988 11200
rect 2380 10388 2436 11200
rect 2380 10332 2548 10388
rect 2150 10220 2414 10230
rect 2206 10164 2254 10220
rect 2310 10164 2358 10220
rect 2150 10154 2414 10164
rect 2150 8652 2414 8662
rect 2206 8596 2254 8652
rect 2310 8596 2358 8652
rect 2150 8586 2414 8596
rect 1932 8318 1934 8370
rect 1986 8318 1988 8370
rect 1932 8306 1988 8318
rect 2150 7084 2414 7094
rect 2206 7028 2254 7084
rect 2310 7028 2358 7084
rect 2150 7018 2414 7028
rect 2492 6802 2548 10332
rect 2828 8930 2884 11200
rect 3276 10052 3332 11200
rect 2828 8878 2830 8930
rect 2882 8878 2884 8930
rect 2828 8866 2884 8878
rect 3052 9996 3332 10052
rect 2828 8708 2884 8718
rect 2716 8148 2772 8158
rect 2604 7364 2660 7374
rect 2604 7270 2660 7308
rect 2492 6750 2494 6802
rect 2546 6750 2548 6802
rect 2492 6738 2548 6750
rect 2604 6692 2660 6702
rect 588 3602 644 3612
rect 1484 3948 1652 4004
rect 1932 6580 1988 6590
rect 1260 3556 1316 3566
rect 700 3554 1316 3556
rect 700 3502 1262 3554
rect 1314 3502 1316 3554
rect 700 3500 1316 3502
rect 700 3444 756 3500
rect 1260 3490 1316 3500
rect 588 3442 756 3444
rect 588 3390 702 3442
rect 754 3390 756 3442
rect 588 3388 756 3390
rect 588 800 644 3388
rect 700 3378 756 3388
rect 812 1988 868 1998
rect 1260 1988 1316 1998
rect 812 1986 1316 1988
rect 812 1934 814 1986
rect 866 1934 1262 1986
rect 1314 1934 1316 1986
rect 812 1932 1316 1934
rect 812 1922 868 1932
rect 1036 800 1092 1932
rect 1260 1922 1316 1932
rect 1484 800 1540 3948
rect 1596 2996 1652 3006
rect 1596 2902 1652 2940
rect 1932 800 1988 6524
rect 2150 5516 2414 5526
rect 2206 5460 2254 5516
rect 2310 5460 2358 5516
rect 2150 5450 2414 5460
rect 2492 5012 2548 5022
rect 2150 3948 2414 3958
rect 2206 3892 2254 3948
rect 2310 3892 2358 3948
rect 2150 3882 2414 3892
rect 2380 3668 2436 3678
rect 2380 3574 2436 3612
rect 2156 2996 2212 3006
rect 2156 2770 2212 2940
rect 2156 2718 2158 2770
rect 2210 2718 2212 2770
rect 2156 2706 2212 2718
rect 2150 2380 2414 2390
rect 2206 2324 2254 2380
rect 2310 2324 2358 2380
rect 2150 2314 2414 2324
rect 2492 2098 2548 4956
rect 2492 2046 2494 2098
rect 2546 2046 2548 2098
rect 2492 2034 2548 2046
rect 2604 1876 2660 6636
rect 2716 5234 2772 8092
rect 2716 5182 2718 5234
rect 2770 5182 2772 5234
rect 2716 5170 2772 5182
rect 2380 1820 2660 1876
rect 2380 800 2436 1820
rect 2828 800 2884 8652
rect 3052 5794 3108 9996
rect 3388 9828 3444 9838
rect 3388 9734 3444 9772
rect 3724 8428 3780 11200
rect 4172 9828 4228 11200
rect 3612 8372 3780 8428
rect 4060 9772 4228 9828
rect 4620 9828 4676 11200
rect 4956 9828 5012 9838
rect 4620 9772 4788 9828
rect 3500 8258 3556 8270
rect 3500 8206 3502 8258
rect 3554 8206 3556 8258
rect 3500 8036 3556 8206
rect 3388 6692 3444 6702
rect 3388 6598 3444 6636
rect 3500 6580 3556 7980
rect 3500 6514 3556 6524
rect 3052 5742 3054 5794
rect 3106 5742 3108 5794
rect 3052 5730 3108 5742
rect 3164 5908 3220 5918
rect 3164 3220 3220 5852
rect 3612 4452 3668 8372
rect 3724 7474 3780 7486
rect 3724 7422 3726 7474
rect 3778 7422 3780 7474
rect 3724 6468 3780 7422
rect 4060 7364 4116 9772
rect 4620 9602 4676 9614
rect 4620 9550 4622 9602
rect 4674 9550 4676 9602
rect 4208 9436 4472 9446
rect 4264 9380 4312 9436
rect 4368 9380 4416 9436
rect 4208 9370 4472 9380
rect 4396 9044 4452 9054
rect 4620 9044 4676 9550
rect 4396 9042 4676 9044
rect 4396 8990 4398 9042
rect 4450 8990 4676 9042
rect 4396 8988 4676 8990
rect 4396 8708 4452 8988
rect 4396 8642 4452 8652
rect 4508 8036 4564 8074
rect 4508 7970 4564 7980
rect 4208 7868 4472 7878
rect 4264 7812 4312 7868
rect 4368 7812 4416 7868
rect 4208 7802 4472 7812
rect 4060 7298 4116 7308
rect 4508 6468 4564 6478
rect 3724 6466 4564 6468
rect 3724 6414 4510 6466
rect 4562 6414 4564 6466
rect 3724 6412 4564 6414
rect 3836 5124 3892 5134
rect 3836 5030 3892 5068
rect 3612 4386 3668 4396
rect 3276 4338 3332 4350
rect 3276 4286 3278 4338
rect 3330 4286 3332 4338
rect 3276 3444 3332 4286
rect 3276 3378 3332 3388
rect 3724 3444 3780 3454
rect 3164 3164 3332 3220
rect 3276 800 3332 3164
rect 3724 800 3780 3388
rect 4060 1428 4116 6412
rect 4508 6402 4564 6412
rect 4208 6300 4472 6310
rect 4264 6244 4312 6300
rect 4368 6244 4416 6300
rect 4208 6234 4472 6244
rect 4172 5908 4228 5918
rect 4172 5814 4228 5852
rect 4508 5124 4564 5134
rect 4508 5030 4564 5068
rect 4208 4732 4472 4742
rect 4264 4676 4312 4732
rect 4368 4676 4416 4732
rect 4208 4666 4472 4676
rect 4620 4340 4676 4350
rect 4508 3444 4564 3454
rect 4508 3350 4564 3388
rect 4208 3164 4472 3174
rect 4264 3108 4312 3164
rect 4368 3108 4416 3164
rect 4208 3098 4472 3108
rect 4508 2660 4564 2670
rect 4508 2566 4564 2604
rect 4208 1596 4472 1606
rect 4264 1540 4312 1596
rect 4368 1540 4416 1596
rect 4208 1530 4472 1540
rect 4060 1372 4228 1428
rect 4172 800 4228 1372
rect 4620 800 4676 4284
rect 4732 4226 4788 9772
rect 5068 9828 5124 11200
rect 5068 9772 5236 9828
rect 4956 9604 5012 9772
rect 5068 9604 5124 9614
rect 4956 9602 5124 9604
rect 4956 9550 5070 9602
rect 5122 9550 5124 9602
rect 4956 9548 5124 9550
rect 5068 9538 5124 9548
rect 5068 8932 5124 8942
rect 5068 8370 5124 8876
rect 5068 8318 5070 8370
rect 5122 8318 5124 8370
rect 5068 8306 5124 8318
rect 5068 7476 5124 7486
rect 4956 6466 5012 6478
rect 4956 6414 4958 6466
rect 5010 6414 5012 6466
rect 4956 5908 5012 6414
rect 4956 5842 5012 5852
rect 4732 4174 4734 4226
rect 4786 4174 4788 4226
rect 4732 4162 4788 4174
rect 5068 800 5124 7420
rect 5180 7362 5236 9772
rect 5292 9042 5348 9054
rect 5292 8990 5294 9042
rect 5346 8990 5348 9042
rect 5292 8932 5348 8990
rect 5292 8866 5348 8876
rect 5180 7310 5182 7362
rect 5234 7310 5236 7362
rect 5180 7298 5236 7310
rect 5404 6692 5460 6702
rect 5404 6598 5460 6636
rect 5516 2098 5572 11200
rect 5964 5234 6020 11200
rect 6412 10388 6468 11200
rect 6076 10332 6468 10388
rect 6076 8148 6132 10332
rect 6266 10220 6530 10230
rect 6322 10164 6370 10220
rect 6426 10164 6474 10220
rect 6266 10154 6530 10164
rect 6266 8652 6530 8662
rect 6322 8596 6370 8652
rect 6426 8596 6474 8652
rect 6266 8586 6530 8596
rect 6860 8428 6916 11200
rect 6076 8082 6132 8092
rect 6636 8372 6916 8428
rect 5964 5182 5966 5234
rect 6018 5182 6020 5234
rect 5964 5170 6020 5182
rect 6076 7588 6132 7598
rect 5964 4788 6020 4798
rect 5852 4340 5908 4350
rect 5852 4246 5908 4284
rect 5516 2046 5518 2098
rect 5570 2046 5572 2098
rect 5516 2034 5572 2046
rect 5516 1876 5572 1886
rect 5516 800 5572 1820
rect 5964 800 6020 4732
rect 6076 2882 6132 7532
rect 6300 7476 6356 7486
rect 6300 7382 6356 7420
rect 6266 7084 6530 7094
rect 6322 7028 6370 7084
rect 6426 7028 6474 7084
rect 6266 7018 6530 7028
rect 6636 5794 6692 8372
rect 7308 7588 7364 11200
rect 7644 8930 7700 8942
rect 7644 8878 7646 8930
rect 7698 8878 7700 8930
rect 7644 8820 7700 8878
rect 7644 8754 7700 8764
rect 7756 8370 7812 11200
rect 7756 8318 7758 8370
rect 7810 8318 7812 8370
rect 7756 8306 7812 8318
rect 7308 7522 7364 7532
rect 7308 7364 7364 7374
rect 7308 7270 7364 7308
rect 8204 6802 8260 11200
rect 8324 9436 8588 9446
rect 8380 9380 8428 9436
rect 8484 9380 8532 9436
rect 8324 9370 8588 9380
rect 8324 7868 8588 7878
rect 8380 7812 8428 7868
rect 8484 7812 8532 7868
rect 8324 7802 8588 7812
rect 8652 6916 8708 11200
rect 8652 6850 8708 6860
rect 8876 8258 8932 8270
rect 8876 8206 8878 8258
rect 8930 8206 8932 8258
rect 8204 6750 8206 6802
rect 8258 6750 8260 6802
rect 8204 6738 8260 6750
rect 7980 6692 8036 6702
rect 6636 5742 6638 5794
rect 6690 5742 6692 5794
rect 6636 5730 6692 5742
rect 7532 5906 7588 5918
rect 7532 5854 7534 5906
rect 7586 5854 7588 5906
rect 6266 5516 6530 5526
rect 6322 5460 6370 5516
rect 6426 5460 6474 5516
rect 6266 5450 6530 5460
rect 6636 5124 6692 5134
rect 6266 3948 6530 3958
rect 6322 3892 6370 3948
rect 6426 3892 6474 3948
rect 6266 3882 6530 3892
rect 6524 3668 6580 3678
rect 6524 3574 6580 3612
rect 6076 2830 6078 2882
rect 6130 2830 6132 2882
rect 6076 2818 6132 2830
rect 6266 2380 6530 2390
rect 6322 2324 6370 2380
rect 6426 2324 6474 2380
rect 6266 2314 6530 2324
rect 6636 2212 6692 5068
rect 7196 5122 7252 5134
rect 7196 5070 7198 5122
rect 7250 5070 7252 5122
rect 7196 4788 7252 5070
rect 7196 4722 7252 4732
rect 6860 4340 6916 4350
rect 6860 4246 6916 4284
rect 6412 2156 6692 2212
rect 6860 4116 6916 4126
rect 6412 800 6468 2156
rect 6748 1986 6804 1998
rect 6748 1934 6750 1986
rect 6802 1934 6804 1986
rect 6748 1876 6804 1934
rect 6748 1810 6804 1820
rect 6860 800 6916 4060
rect 7532 4116 7588 5854
rect 7868 4564 7924 4574
rect 7532 4050 7588 4060
rect 7644 4508 7868 4564
rect 7644 3554 7700 4508
rect 7868 4470 7924 4508
rect 7644 3502 7646 3554
rect 7698 3502 7700 3554
rect 7644 3490 7700 3502
rect 7308 2772 7364 2782
rect 7308 800 7364 2716
rect 7756 1876 7812 1886
rect 7756 1782 7812 1820
rect 7980 1652 8036 6636
rect 8876 6692 8932 8206
rect 8876 6626 8932 6636
rect 7756 1596 8036 1652
rect 8204 6580 8260 6590
rect 7756 800 7812 1596
rect 8204 800 8260 6524
rect 8324 6300 8588 6310
rect 8380 6244 8428 6300
rect 8484 6244 8532 6300
rect 8324 6234 8588 6244
rect 8988 4900 9044 4910
rect 8324 4732 8588 4742
rect 8380 4676 8428 4732
rect 8484 4676 8532 4732
rect 8324 4666 8588 4676
rect 8988 4562 9044 4844
rect 8988 4510 8990 4562
rect 9042 4510 9044 4562
rect 8988 4498 9044 4510
rect 8540 4226 8596 4238
rect 8540 4174 8542 4226
rect 8594 4174 8596 4226
rect 8540 4116 8596 4174
rect 9100 4228 9156 11200
rect 9548 6804 9604 11200
rect 9548 6738 9604 6748
rect 9884 8034 9940 8046
rect 9884 7982 9886 8034
rect 9938 7982 9940 8034
rect 9324 6690 9380 6702
rect 9324 6638 9326 6690
rect 9378 6638 9380 6690
rect 9324 6580 9380 6638
rect 9884 6692 9940 7982
rect 9884 6626 9940 6636
rect 9324 6514 9380 6524
rect 9996 6468 10052 11200
rect 10444 10388 10500 11200
rect 9996 6402 10052 6412
rect 10220 10332 10500 10388
rect 9996 5794 10052 5806
rect 9996 5742 9998 5794
rect 10050 5742 10052 5794
rect 9100 4162 9156 4172
rect 9548 5234 9604 5246
rect 9548 5182 9550 5234
rect 9602 5182 9604 5234
rect 8540 4050 8596 4060
rect 9100 3666 9156 3678
rect 9100 3614 9102 3666
rect 9154 3614 9156 3666
rect 8324 3164 8588 3174
rect 8380 3108 8428 3164
rect 8484 3108 8532 3164
rect 8324 3098 8588 3108
rect 8540 2772 8596 2782
rect 8540 2678 8596 2716
rect 8764 2100 8820 2110
rect 8652 2098 8820 2100
rect 8652 2046 8766 2098
rect 8818 2046 8820 2098
rect 8652 2044 8820 2046
rect 8324 1596 8588 1606
rect 8380 1540 8428 1596
rect 8484 1540 8532 1596
rect 8324 1530 8588 1540
rect 8652 800 8708 2044
rect 8764 2034 8820 2044
rect 9100 800 9156 3614
rect 9548 800 9604 5182
rect 9996 800 10052 5742
rect 10220 4564 10276 10332
rect 10382 10220 10646 10230
rect 10438 10164 10486 10220
rect 10542 10164 10590 10220
rect 10382 10154 10646 10164
rect 10780 8930 10836 8942
rect 10780 8878 10782 8930
rect 10834 8878 10836 8930
rect 10382 8652 10646 8662
rect 10438 8596 10486 8652
rect 10542 8596 10590 8652
rect 10382 8586 10646 8596
rect 10780 8484 10836 8878
rect 10780 8418 10836 8428
rect 10382 7084 10646 7094
rect 10438 7028 10486 7084
rect 10542 7028 10590 7084
rect 10382 7018 10646 7028
rect 10892 7028 10948 11200
rect 11340 9380 11396 11200
rect 11788 9828 11844 11200
rect 11788 9772 12068 9828
rect 11676 9716 11732 9726
rect 11340 9324 11508 9380
rect 11452 8428 11508 9324
rect 11676 9044 11732 9660
rect 11676 9042 11956 9044
rect 11676 8990 11678 9042
rect 11730 8990 11956 9042
rect 11676 8988 11956 8990
rect 11676 8978 11732 8988
rect 11452 8372 11844 8428
rect 10892 6962 10948 6972
rect 11676 7028 11732 7038
rect 11116 6916 11172 6926
rect 10780 6804 10836 6814
rect 10332 6580 10388 6590
rect 10332 6486 10388 6524
rect 10382 5516 10646 5526
rect 10438 5460 10486 5516
rect 10542 5460 10590 5516
rect 10382 5450 10646 5460
rect 10220 4498 10276 4508
rect 10780 5122 10836 6748
rect 11004 6468 11060 6478
rect 11004 5906 11060 6412
rect 11004 5854 11006 5906
rect 11058 5854 11060 5906
rect 11004 5236 11060 5854
rect 11004 5170 11060 5180
rect 10780 5070 10782 5122
rect 10834 5070 10836 5122
rect 10220 4228 10276 4238
rect 10108 3668 10164 3678
rect 10108 1876 10164 3612
rect 10220 3556 10276 4172
rect 10382 3948 10646 3958
rect 10438 3892 10486 3948
rect 10542 3892 10590 3948
rect 10382 3882 10646 3892
rect 10780 3666 10836 5070
rect 10780 3614 10782 3666
rect 10834 3614 10836 3666
rect 10780 3602 10836 3614
rect 10220 3424 10276 3500
rect 10892 2658 10948 2670
rect 10892 2606 10894 2658
rect 10946 2606 10948 2658
rect 10382 2380 10646 2390
rect 10438 2324 10486 2380
rect 10542 2324 10590 2380
rect 10382 2314 10646 2324
rect 10108 1820 10500 1876
rect 10444 800 10500 1820
rect 10892 800 10948 2606
rect 11116 2098 11172 6860
rect 11452 4564 11508 4574
rect 11228 3668 11284 3678
rect 11228 3666 11396 3668
rect 11228 3614 11230 3666
rect 11282 3614 11396 3666
rect 11228 3612 11396 3614
rect 11228 3602 11284 3612
rect 11340 3554 11396 3612
rect 11340 3502 11342 3554
rect 11394 3502 11396 3554
rect 11340 3490 11396 3502
rect 11452 2884 11508 4508
rect 11676 3332 11732 6972
rect 11788 6804 11844 8372
rect 11900 8370 11956 8988
rect 11900 8318 11902 8370
rect 11954 8318 11956 8370
rect 11900 8306 11956 8318
rect 11788 6690 11844 6748
rect 11788 6638 11790 6690
rect 11842 6638 11844 6690
rect 11788 6626 11844 6638
rect 11788 5236 11844 5246
rect 11788 5142 11844 5180
rect 12012 4340 12068 9772
rect 12236 7700 12292 11200
rect 12684 9828 12740 11200
rect 12684 9772 12852 9828
rect 12440 9436 12704 9446
rect 12496 9380 12544 9436
rect 12600 9380 12648 9436
rect 12440 9370 12704 9380
rect 12796 8260 12852 9772
rect 13132 8428 13188 11200
rect 13132 8372 13300 8428
rect 12796 8194 12852 8204
rect 12440 7868 12704 7878
rect 12496 7812 12544 7868
rect 12600 7812 12648 7868
rect 12440 7802 12704 7812
rect 12236 7634 12292 7644
rect 13132 7700 13188 7710
rect 13132 7474 13188 7644
rect 13132 7422 13134 7474
rect 13186 7422 13188 7474
rect 13132 7410 13188 7422
rect 12236 7362 12292 7374
rect 12236 7310 12238 7362
rect 12290 7310 12292 7362
rect 12124 6804 12180 6814
rect 12124 5906 12180 6748
rect 12124 5854 12126 5906
rect 12178 5854 12180 5906
rect 12124 5842 12180 5854
rect 12012 4274 12068 4284
rect 11900 4226 11956 4238
rect 11900 4174 11902 4226
rect 11954 4174 11956 4226
rect 11788 3556 11844 3566
rect 11788 3462 11844 3500
rect 11788 3332 11844 3342
rect 11676 3276 11788 3332
rect 11788 3266 11844 3276
rect 11900 2996 11956 4174
rect 11116 2046 11118 2098
rect 11170 2046 11172 2098
rect 11116 1986 11172 2046
rect 11116 1934 11118 1986
rect 11170 1934 11172 1986
rect 11116 1922 11172 1934
rect 11340 2828 11508 2884
rect 11788 2940 11956 2996
rect 12012 3332 12068 3342
rect 11340 800 11396 2828
rect 11452 2100 11508 2110
rect 11452 2098 11620 2100
rect 11452 2046 11454 2098
rect 11506 2046 11620 2098
rect 11452 2044 11620 2046
rect 11452 2034 11508 2044
rect 11564 1986 11620 2044
rect 11564 1934 11566 1986
rect 11618 1934 11620 1986
rect 11564 1922 11620 1934
rect 11788 800 11844 2940
rect 12012 2770 12068 3276
rect 12012 2718 12014 2770
rect 12066 2718 12068 2770
rect 12012 2706 12068 2718
rect 12236 800 12292 7310
rect 13132 6802 13188 6814
rect 13132 6750 13134 6802
rect 13186 6750 13188 6802
rect 12440 6300 12704 6310
rect 12496 6244 12544 6300
rect 12600 6244 12648 6300
rect 12440 6234 12704 6244
rect 12796 5124 12852 5134
rect 12440 4732 12704 4742
rect 12496 4676 12544 4732
rect 12600 4676 12648 4732
rect 12440 4666 12704 4676
rect 12684 4340 12740 4350
rect 12684 4246 12740 4284
rect 12440 3164 12704 3174
rect 12496 3108 12544 3164
rect 12600 3108 12648 3164
rect 12440 3098 12704 3108
rect 12440 1596 12704 1606
rect 12496 1540 12544 1596
rect 12600 1540 12648 1596
rect 12440 1530 12704 1540
rect 12796 1428 12852 5068
rect 12684 1372 12852 1428
rect 12684 800 12740 1372
rect 13132 800 13188 6750
rect 13244 6692 13300 8372
rect 13244 6626 13300 6636
rect 13468 8370 13524 8382
rect 13468 8318 13470 8370
rect 13522 8318 13524 8370
rect 13468 5124 13524 8318
rect 13468 5058 13524 5068
rect 13580 4116 13636 11200
rect 13916 9938 13972 9950
rect 13916 9886 13918 9938
rect 13970 9886 13972 9938
rect 13916 9156 13972 9886
rect 13916 9090 13972 9100
rect 13916 8930 13972 8942
rect 13916 8878 13918 8930
rect 13970 8878 13972 8930
rect 13916 6020 13972 8878
rect 14028 6244 14084 11200
rect 14476 10388 14532 11200
rect 14364 10332 14532 10388
rect 14364 9044 14420 10332
rect 14498 10220 14762 10230
rect 14554 10164 14602 10220
rect 14658 10164 14706 10220
rect 14498 10154 14762 10164
rect 14924 9940 14980 11200
rect 14924 9826 14980 9884
rect 14924 9774 14926 9826
rect 14978 9774 14980 9826
rect 14924 9762 14980 9774
rect 14924 9156 14980 9166
rect 14476 9044 14532 9054
rect 14364 8988 14476 9044
rect 14476 8912 14532 8988
rect 14498 8652 14762 8662
rect 14554 8596 14602 8652
rect 14658 8596 14706 8652
rect 14498 8586 14762 8596
rect 14588 8260 14644 8270
rect 14588 8166 14644 8204
rect 14140 7700 14196 7710
rect 14140 7606 14196 7644
rect 14498 7084 14762 7094
rect 14554 7028 14602 7084
rect 14658 7028 14706 7084
rect 14498 7018 14762 7028
rect 14588 6692 14644 6702
rect 14588 6598 14644 6636
rect 14028 6178 14084 6188
rect 13916 5964 14420 6020
rect 13692 5794 13748 5806
rect 13692 5742 13694 5794
rect 13746 5742 13748 5794
rect 13692 4564 13748 5742
rect 13692 4498 13748 4508
rect 14028 5234 14084 5246
rect 14028 5182 14030 5234
rect 14082 5182 14084 5234
rect 13692 4340 13748 4350
rect 13692 4246 13748 4284
rect 13580 4060 13748 4116
rect 13580 3666 13636 3678
rect 13580 3614 13582 3666
rect 13634 3614 13636 3666
rect 13580 800 13636 3614
rect 13692 3556 13748 4060
rect 13692 3490 13748 3500
rect 13916 2100 13972 2110
rect 13916 2006 13972 2044
rect 14028 800 14084 5182
rect 14140 4226 14196 4238
rect 14140 4174 14142 4226
rect 14194 4174 14196 4226
rect 14140 3332 14196 4174
rect 14140 3266 14196 3276
rect 14364 1764 14420 5964
rect 14498 5516 14762 5526
rect 14554 5460 14602 5516
rect 14658 5460 14706 5516
rect 14498 5450 14762 5460
rect 14498 3948 14762 3958
rect 14554 3892 14602 3948
rect 14658 3892 14706 3948
rect 14498 3882 14762 3892
rect 14588 3556 14644 3566
rect 14588 3462 14644 3500
rect 14476 2660 14532 2670
rect 14476 2566 14532 2604
rect 14498 2380 14762 2390
rect 14554 2324 14602 2380
rect 14658 2324 14706 2380
rect 14498 2314 14762 2324
rect 14364 1708 14532 1764
rect 14476 800 14532 1708
rect 14924 800 14980 9100
rect 15036 6244 15092 6254
rect 15036 5236 15092 6188
rect 15036 5122 15092 5180
rect 15036 5070 15038 5122
rect 15090 5070 15092 5122
rect 15036 5058 15092 5070
rect 15372 3780 15428 11200
rect 15484 9940 15540 9950
rect 15484 9846 15540 9884
rect 15484 9044 15540 9054
rect 15484 8950 15540 8988
rect 15820 8428 15876 11200
rect 16268 9716 16324 11200
rect 16268 9650 16324 9660
rect 16556 9436 16820 9446
rect 16612 9380 16660 9436
rect 16716 9380 16764 9436
rect 16556 9370 16820 9380
rect 15708 8372 15876 8428
rect 16156 8484 16212 8494
rect 16156 8372 16324 8428
rect 15596 8260 15652 8270
rect 15596 8166 15652 8204
rect 15596 6692 15652 6702
rect 15596 6598 15652 6636
rect 15596 5236 15652 5246
rect 15596 5142 15652 5180
rect 15372 3778 15540 3780
rect 15372 3726 15374 3778
rect 15426 3726 15540 3778
rect 15372 3724 15540 3726
rect 15372 3714 15428 3724
rect 15484 2770 15540 3724
rect 15596 3556 15652 3566
rect 15596 3462 15652 3500
rect 15484 2718 15486 2770
rect 15538 2718 15540 2770
rect 15484 2706 15540 2718
rect 15372 2660 15428 2670
rect 15036 1988 15092 1998
rect 15036 1894 15092 1932
rect 15372 800 15428 2604
rect 15596 2100 15652 2110
rect 15708 2100 15764 8372
rect 16044 3778 16100 3790
rect 16044 3726 16046 3778
rect 16098 3726 16100 3778
rect 16044 3666 16100 3726
rect 16044 3614 16046 3666
rect 16098 3614 16100 3666
rect 16044 3602 16100 3614
rect 15596 2098 15764 2100
rect 15596 2046 15598 2098
rect 15650 2046 15764 2098
rect 15596 2044 15764 2046
rect 15820 2100 15876 2110
rect 15596 1988 15652 2044
rect 15596 1922 15652 1932
rect 15820 800 15876 2044
rect 16268 800 16324 8372
rect 16556 7868 16820 7878
rect 16612 7812 16660 7868
rect 16716 7812 16764 7868
rect 16556 7802 16820 7812
rect 16556 6300 16820 6310
rect 16612 6244 16660 6300
rect 16716 6244 16764 6300
rect 16556 6234 16820 6244
rect 16556 4732 16820 4742
rect 16612 4676 16660 4732
rect 16716 4676 16764 4732
rect 16556 4666 16820 4676
rect 16556 3164 16820 3174
rect 16612 3108 16660 3164
rect 16716 3108 16764 3164
rect 16556 3098 16820 3108
rect 16556 1596 16820 1606
rect 16612 1540 16660 1596
rect 16716 1540 16764 1596
rect 16556 1530 16820 1540
rect 560 0 672 800
rect 1008 0 1120 800
rect 1456 0 1568 800
rect 1904 0 2016 800
rect 2352 0 2464 800
rect 2800 0 2912 800
rect 3248 0 3360 800
rect 3696 0 3808 800
rect 4144 0 4256 800
rect 4592 0 4704 800
rect 5040 0 5152 800
rect 5488 0 5600 800
rect 5936 0 6048 800
rect 6384 0 6496 800
rect 6832 0 6944 800
rect 7280 0 7392 800
rect 7728 0 7840 800
rect 8176 0 8288 800
rect 8624 0 8736 800
rect 9072 0 9184 800
rect 9520 0 9632 800
rect 9968 0 10080 800
rect 10416 0 10528 800
rect 10864 0 10976 800
rect 11312 0 11424 800
rect 11760 0 11872 800
rect 12208 0 12320 800
rect 12656 0 12768 800
rect 13104 0 13216 800
rect 13552 0 13664 800
rect 14000 0 14112 800
rect 14448 0 14560 800
rect 14896 0 15008 800
rect 15344 0 15456 800
rect 15792 0 15904 800
rect 16240 0 16352 800
<< via2 >>
rect 1036 4956 1092 5012
rect 1596 9772 1652 9828
rect 1484 4450 1540 4452
rect 1484 4398 1486 4450
rect 1486 4398 1538 4450
rect 1538 4398 1540 4450
rect 1484 4396 1540 4398
rect 2150 10218 2206 10220
rect 2150 10166 2152 10218
rect 2152 10166 2204 10218
rect 2204 10166 2206 10218
rect 2150 10164 2206 10166
rect 2254 10218 2310 10220
rect 2254 10166 2256 10218
rect 2256 10166 2308 10218
rect 2308 10166 2310 10218
rect 2254 10164 2310 10166
rect 2358 10218 2414 10220
rect 2358 10166 2360 10218
rect 2360 10166 2412 10218
rect 2412 10166 2414 10218
rect 2358 10164 2414 10166
rect 2150 8650 2206 8652
rect 2150 8598 2152 8650
rect 2152 8598 2204 8650
rect 2204 8598 2206 8650
rect 2150 8596 2206 8598
rect 2254 8650 2310 8652
rect 2254 8598 2256 8650
rect 2256 8598 2308 8650
rect 2308 8598 2310 8650
rect 2254 8596 2310 8598
rect 2358 8650 2414 8652
rect 2358 8598 2360 8650
rect 2360 8598 2412 8650
rect 2412 8598 2414 8650
rect 2358 8596 2414 8598
rect 2150 7082 2206 7084
rect 2150 7030 2152 7082
rect 2152 7030 2204 7082
rect 2204 7030 2206 7082
rect 2150 7028 2206 7030
rect 2254 7082 2310 7084
rect 2254 7030 2256 7082
rect 2256 7030 2308 7082
rect 2308 7030 2310 7082
rect 2254 7028 2310 7030
rect 2358 7082 2414 7084
rect 2358 7030 2360 7082
rect 2360 7030 2412 7082
rect 2412 7030 2414 7082
rect 2358 7028 2414 7030
rect 2828 8652 2884 8708
rect 2716 8092 2772 8148
rect 2604 7362 2660 7364
rect 2604 7310 2606 7362
rect 2606 7310 2658 7362
rect 2658 7310 2660 7362
rect 2604 7308 2660 7310
rect 2604 6636 2660 6692
rect 588 3612 644 3668
rect 1932 6524 1988 6580
rect 1596 2994 1652 2996
rect 1596 2942 1598 2994
rect 1598 2942 1650 2994
rect 1650 2942 1652 2994
rect 1596 2940 1652 2942
rect 2150 5514 2206 5516
rect 2150 5462 2152 5514
rect 2152 5462 2204 5514
rect 2204 5462 2206 5514
rect 2150 5460 2206 5462
rect 2254 5514 2310 5516
rect 2254 5462 2256 5514
rect 2256 5462 2308 5514
rect 2308 5462 2310 5514
rect 2254 5460 2310 5462
rect 2358 5514 2414 5516
rect 2358 5462 2360 5514
rect 2360 5462 2412 5514
rect 2412 5462 2414 5514
rect 2358 5460 2414 5462
rect 2492 4956 2548 5012
rect 2150 3946 2206 3948
rect 2150 3894 2152 3946
rect 2152 3894 2204 3946
rect 2204 3894 2206 3946
rect 2150 3892 2206 3894
rect 2254 3946 2310 3948
rect 2254 3894 2256 3946
rect 2256 3894 2308 3946
rect 2308 3894 2310 3946
rect 2254 3892 2310 3894
rect 2358 3946 2414 3948
rect 2358 3894 2360 3946
rect 2360 3894 2412 3946
rect 2412 3894 2414 3946
rect 2358 3892 2414 3894
rect 2380 3666 2436 3668
rect 2380 3614 2382 3666
rect 2382 3614 2434 3666
rect 2434 3614 2436 3666
rect 2380 3612 2436 3614
rect 2156 2940 2212 2996
rect 2150 2378 2206 2380
rect 2150 2326 2152 2378
rect 2152 2326 2204 2378
rect 2204 2326 2206 2378
rect 2150 2324 2206 2326
rect 2254 2378 2310 2380
rect 2254 2326 2256 2378
rect 2256 2326 2308 2378
rect 2308 2326 2310 2378
rect 2254 2324 2310 2326
rect 2358 2378 2414 2380
rect 2358 2326 2360 2378
rect 2360 2326 2412 2378
rect 2412 2326 2414 2378
rect 2358 2324 2414 2326
rect 3388 9826 3444 9828
rect 3388 9774 3390 9826
rect 3390 9774 3442 9826
rect 3442 9774 3444 9826
rect 3388 9772 3444 9774
rect 3500 7980 3556 8036
rect 3388 6690 3444 6692
rect 3388 6638 3390 6690
rect 3390 6638 3442 6690
rect 3442 6638 3444 6690
rect 3388 6636 3444 6638
rect 3500 6524 3556 6580
rect 3164 5852 3220 5908
rect 4208 9434 4264 9436
rect 4208 9382 4210 9434
rect 4210 9382 4262 9434
rect 4262 9382 4264 9434
rect 4208 9380 4264 9382
rect 4312 9434 4368 9436
rect 4312 9382 4314 9434
rect 4314 9382 4366 9434
rect 4366 9382 4368 9434
rect 4312 9380 4368 9382
rect 4416 9434 4472 9436
rect 4416 9382 4418 9434
rect 4418 9382 4470 9434
rect 4470 9382 4472 9434
rect 4416 9380 4472 9382
rect 4396 8652 4452 8708
rect 4508 8034 4564 8036
rect 4508 7982 4510 8034
rect 4510 7982 4562 8034
rect 4562 7982 4564 8034
rect 4508 7980 4564 7982
rect 4208 7866 4264 7868
rect 4208 7814 4210 7866
rect 4210 7814 4262 7866
rect 4262 7814 4264 7866
rect 4208 7812 4264 7814
rect 4312 7866 4368 7868
rect 4312 7814 4314 7866
rect 4314 7814 4366 7866
rect 4366 7814 4368 7866
rect 4312 7812 4368 7814
rect 4416 7866 4472 7868
rect 4416 7814 4418 7866
rect 4418 7814 4470 7866
rect 4470 7814 4472 7866
rect 4416 7812 4472 7814
rect 4060 7308 4116 7364
rect 3836 5122 3892 5124
rect 3836 5070 3838 5122
rect 3838 5070 3890 5122
rect 3890 5070 3892 5122
rect 3836 5068 3892 5070
rect 3612 4396 3668 4452
rect 3276 3388 3332 3444
rect 3724 3388 3780 3444
rect 4208 6298 4264 6300
rect 4208 6246 4210 6298
rect 4210 6246 4262 6298
rect 4262 6246 4264 6298
rect 4208 6244 4264 6246
rect 4312 6298 4368 6300
rect 4312 6246 4314 6298
rect 4314 6246 4366 6298
rect 4366 6246 4368 6298
rect 4312 6244 4368 6246
rect 4416 6298 4472 6300
rect 4416 6246 4418 6298
rect 4418 6246 4470 6298
rect 4470 6246 4472 6298
rect 4416 6244 4472 6246
rect 4172 5906 4228 5908
rect 4172 5854 4174 5906
rect 4174 5854 4226 5906
rect 4226 5854 4228 5906
rect 4172 5852 4228 5854
rect 4508 5122 4564 5124
rect 4508 5070 4510 5122
rect 4510 5070 4562 5122
rect 4562 5070 4564 5122
rect 4508 5068 4564 5070
rect 4208 4730 4264 4732
rect 4208 4678 4210 4730
rect 4210 4678 4262 4730
rect 4262 4678 4264 4730
rect 4208 4676 4264 4678
rect 4312 4730 4368 4732
rect 4312 4678 4314 4730
rect 4314 4678 4366 4730
rect 4366 4678 4368 4730
rect 4312 4676 4368 4678
rect 4416 4730 4472 4732
rect 4416 4678 4418 4730
rect 4418 4678 4470 4730
rect 4470 4678 4472 4730
rect 4416 4676 4472 4678
rect 4620 4284 4676 4340
rect 4508 3442 4564 3444
rect 4508 3390 4510 3442
rect 4510 3390 4562 3442
rect 4562 3390 4564 3442
rect 4508 3388 4564 3390
rect 4208 3162 4264 3164
rect 4208 3110 4210 3162
rect 4210 3110 4262 3162
rect 4262 3110 4264 3162
rect 4208 3108 4264 3110
rect 4312 3162 4368 3164
rect 4312 3110 4314 3162
rect 4314 3110 4366 3162
rect 4366 3110 4368 3162
rect 4312 3108 4368 3110
rect 4416 3162 4472 3164
rect 4416 3110 4418 3162
rect 4418 3110 4470 3162
rect 4470 3110 4472 3162
rect 4416 3108 4472 3110
rect 4508 2658 4564 2660
rect 4508 2606 4510 2658
rect 4510 2606 4562 2658
rect 4562 2606 4564 2658
rect 4508 2604 4564 2606
rect 4208 1594 4264 1596
rect 4208 1542 4210 1594
rect 4210 1542 4262 1594
rect 4262 1542 4264 1594
rect 4208 1540 4264 1542
rect 4312 1594 4368 1596
rect 4312 1542 4314 1594
rect 4314 1542 4366 1594
rect 4366 1542 4368 1594
rect 4312 1540 4368 1542
rect 4416 1594 4472 1596
rect 4416 1542 4418 1594
rect 4418 1542 4470 1594
rect 4470 1542 4472 1594
rect 4416 1540 4472 1542
rect 4956 9772 5012 9828
rect 5068 8876 5124 8932
rect 5068 7420 5124 7476
rect 4956 5852 5012 5908
rect 5292 8876 5348 8932
rect 5404 6690 5460 6692
rect 5404 6638 5406 6690
rect 5406 6638 5458 6690
rect 5458 6638 5460 6690
rect 5404 6636 5460 6638
rect 6266 10218 6322 10220
rect 6266 10166 6268 10218
rect 6268 10166 6320 10218
rect 6320 10166 6322 10218
rect 6266 10164 6322 10166
rect 6370 10218 6426 10220
rect 6370 10166 6372 10218
rect 6372 10166 6424 10218
rect 6424 10166 6426 10218
rect 6370 10164 6426 10166
rect 6474 10218 6530 10220
rect 6474 10166 6476 10218
rect 6476 10166 6528 10218
rect 6528 10166 6530 10218
rect 6474 10164 6530 10166
rect 6266 8650 6322 8652
rect 6266 8598 6268 8650
rect 6268 8598 6320 8650
rect 6320 8598 6322 8650
rect 6266 8596 6322 8598
rect 6370 8650 6426 8652
rect 6370 8598 6372 8650
rect 6372 8598 6424 8650
rect 6424 8598 6426 8650
rect 6370 8596 6426 8598
rect 6474 8650 6530 8652
rect 6474 8598 6476 8650
rect 6476 8598 6528 8650
rect 6528 8598 6530 8650
rect 6474 8596 6530 8598
rect 6076 8092 6132 8148
rect 6076 7532 6132 7588
rect 5964 4732 6020 4788
rect 5852 4338 5908 4340
rect 5852 4286 5854 4338
rect 5854 4286 5906 4338
rect 5906 4286 5908 4338
rect 5852 4284 5908 4286
rect 5516 1820 5572 1876
rect 6300 7474 6356 7476
rect 6300 7422 6302 7474
rect 6302 7422 6354 7474
rect 6354 7422 6356 7474
rect 6300 7420 6356 7422
rect 6266 7082 6322 7084
rect 6266 7030 6268 7082
rect 6268 7030 6320 7082
rect 6320 7030 6322 7082
rect 6266 7028 6322 7030
rect 6370 7082 6426 7084
rect 6370 7030 6372 7082
rect 6372 7030 6424 7082
rect 6424 7030 6426 7082
rect 6370 7028 6426 7030
rect 6474 7082 6530 7084
rect 6474 7030 6476 7082
rect 6476 7030 6528 7082
rect 6528 7030 6530 7082
rect 6474 7028 6530 7030
rect 7644 8764 7700 8820
rect 7308 7532 7364 7588
rect 7308 7362 7364 7364
rect 7308 7310 7310 7362
rect 7310 7310 7362 7362
rect 7362 7310 7364 7362
rect 7308 7308 7364 7310
rect 8324 9434 8380 9436
rect 8324 9382 8326 9434
rect 8326 9382 8378 9434
rect 8378 9382 8380 9434
rect 8324 9380 8380 9382
rect 8428 9434 8484 9436
rect 8428 9382 8430 9434
rect 8430 9382 8482 9434
rect 8482 9382 8484 9434
rect 8428 9380 8484 9382
rect 8532 9434 8588 9436
rect 8532 9382 8534 9434
rect 8534 9382 8586 9434
rect 8586 9382 8588 9434
rect 8532 9380 8588 9382
rect 8324 7866 8380 7868
rect 8324 7814 8326 7866
rect 8326 7814 8378 7866
rect 8378 7814 8380 7866
rect 8324 7812 8380 7814
rect 8428 7866 8484 7868
rect 8428 7814 8430 7866
rect 8430 7814 8482 7866
rect 8482 7814 8484 7866
rect 8428 7812 8484 7814
rect 8532 7866 8588 7868
rect 8532 7814 8534 7866
rect 8534 7814 8586 7866
rect 8586 7814 8588 7866
rect 8532 7812 8588 7814
rect 8652 6860 8708 6916
rect 7980 6636 8036 6692
rect 6266 5514 6322 5516
rect 6266 5462 6268 5514
rect 6268 5462 6320 5514
rect 6320 5462 6322 5514
rect 6266 5460 6322 5462
rect 6370 5514 6426 5516
rect 6370 5462 6372 5514
rect 6372 5462 6424 5514
rect 6424 5462 6426 5514
rect 6370 5460 6426 5462
rect 6474 5514 6530 5516
rect 6474 5462 6476 5514
rect 6476 5462 6528 5514
rect 6528 5462 6530 5514
rect 6474 5460 6530 5462
rect 6636 5068 6692 5124
rect 6266 3946 6322 3948
rect 6266 3894 6268 3946
rect 6268 3894 6320 3946
rect 6320 3894 6322 3946
rect 6266 3892 6322 3894
rect 6370 3946 6426 3948
rect 6370 3894 6372 3946
rect 6372 3894 6424 3946
rect 6424 3894 6426 3946
rect 6370 3892 6426 3894
rect 6474 3946 6530 3948
rect 6474 3894 6476 3946
rect 6476 3894 6528 3946
rect 6528 3894 6530 3946
rect 6474 3892 6530 3894
rect 6524 3666 6580 3668
rect 6524 3614 6526 3666
rect 6526 3614 6578 3666
rect 6578 3614 6580 3666
rect 6524 3612 6580 3614
rect 6266 2378 6322 2380
rect 6266 2326 6268 2378
rect 6268 2326 6320 2378
rect 6320 2326 6322 2378
rect 6266 2324 6322 2326
rect 6370 2378 6426 2380
rect 6370 2326 6372 2378
rect 6372 2326 6424 2378
rect 6424 2326 6426 2378
rect 6370 2324 6426 2326
rect 6474 2378 6530 2380
rect 6474 2326 6476 2378
rect 6476 2326 6528 2378
rect 6528 2326 6530 2378
rect 6474 2324 6530 2326
rect 7196 4732 7252 4788
rect 6860 4338 6916 4340
rect 6860 4286 6862 4338
rect 6862 4286 6914 4338
rect 6914 4286 6916 4338
rect 6860 4284 6916 4286
rect 6860 4060 6916 4116
rect 6748 1820 6804 1876
rect 7532 4060 7588 4116
rect 7868 4562 7924 4564
rect 7868 4510 7870 4562
rect 7870 4510 7922 4562
rect 7922 4510 7924 4562
rect 7868 4508 7924 4510
rect 7308 2770 7364 2772
rect 7308 2718 7310 2770
rect 7310 2718 7362 2770
rect 7362 2718 7364 2770
rect 7308 2716 7364 2718
rect 7756 1874 7812 1876
rect 7756 1822 7758 1874
rect 7758 1822 7810 1874
rect 7810 1822 7812 1874
rect 7756 1820 7812 1822
rect 8876 6636 8932 6692
rect 8204 6524 8260 6580
rect 8324 6298 8380 6300
rect 8324 6246 8326 6298
rect 8326 6246 8378 6298
rect 8378 6246 8380 6298
rect 8324 6244 8380 6246
rect 8428 6298 8484 6300
rect 8428 6246 8430 6298
rect 8430 6246 8482 6298
rect 8482 6246 8484 6298
rect 8428 6244 8484 6246
rect 8532 6298 8588 6300
rect 8532 6246 8534 6298
rect 8534 6246 8586 6298
rect 8586 6246 8588 6298
rect 8532 6244 8588 6246
rect 8988 4844 9044 4900
rect 8324 4730 8380 4732
rect 8324 4678 8326 4730
rect 8326 4678 8378 4730
rect 8378 4678 8380 4730
rect 8324 4676 8380 4678
rect 8428 4730 8484 4732
rect 8428 4678 8430 4730
rect 8430 4678 8482 4730
rect 8482 4678 8484 4730
rect 8428 4676 8484 4678
rect 8532 4730 8588 4732
rect 8532 4678 8534 4730
rect 8534 4678 8586 4730
rect 8586 4678 8588 4730
rect 8532 4676 8588 4678
rect 9548 6748 9604 6804
rect 9884 6636 9940 6692
rect 9324 6524 9380 6580
rect 9996 6412 10052 6468
rect 9100 4172 9156 4228
rect 8540 4060 8596 4116
rect 8324 3162 8380 3164
rect 8324 3110 8326 3162
rect 8326 3110 8378 3162
rect 8378 3110 8380 3162
rect 8324 3108 8380 3110
rect 8428 3162 8484 3164
rect 8428 3110 8430 3162
rect 8430 3110 8482 3162
rect 8482 3110 8484 3162
rect 8428 3108 8484 3110
rect 8532 3162 8588 3164
rect 8532 3110 8534 3162
rect 8534 3110 8586 3162
rect 8586 3110 8588 3162
rect 8532 3108 8588 3110
rect 8540 2770 8596 2772
rect 8540 2718 8542 2770
rect 8542 2718 8594 2770
rect 8594 2718 8596 2770
rect 8540 2716 8596 2718
rect 8324 1594 8380 1596
rect 8324 1542 8326 1594
rect 8326 1542 8378 1594
rect 8378 1542 8380 1594
rect 8324 1540 8380 1542
rect 8428 1594 8484 1596
rect 8428 1542 8430 1594
rect 8430 1542 8482 1594
rect 8482 1542 8484 1594
rect 8428 1540 8484 1542
rect 8532 1594 8588 1596
rect 8532 1542 8534 1594
rect 8534 1542 8586 1594
rect 8586 1542 8588 1594
rect 8532 1540 8588 1542
rect 10382 10218 10438 10220
rect 10382 10166 10384 10218
rect 10384 10166 10436 10218
rect 10436 10166 10438 10218
rect 10382 10164 10438 10166
rect 10486 10218 10542 10220
rect 10486 10166 10488 10218
rect 10488 10166 10540 10218
rect 10540 10166 10542 10218
rect 10486 10164 10542 10166
rect 10590 10218 10646 10220
rect 10590 10166 10592 10218
rect 10592 10166 10644 10218
rect 10644 10166 10646 10218
rect 10590 10164 10646 10166
rect 10382 8650 10438 8652
rect 10382 8598 10384 8650
rect 10384 8598 10436 8650
rect 10436 8598 10438 8650
rect 10382 8596 10438 8598
rect 10486 8650 10542 8652
rect 10486 8598 10488 8650
rect 10488 8598 10540 8650
rect 10540 8598 10542 8650
rect 10486 8596 10542 8598
rect 10590 8650 10646 8652
rect 10590 8598 10592 8650
rect 10592 8598 10644 8650
rect 10644 8598 10646 8650
rect 10590 8596 10646 8598
rect 10780 8428 10836 8484
rect 10382 7082 10438 7084
rect 10382 7030 10384 7082
rect 10384 7030 10436 7082
rect 10436 7030 10438 7082
rect 10382 7028 10438 7030
rect 10486 7082 10542 7084
rect 10486 7030 10488 7082
rect 10488 7030 10540 7082
rect 10540 7030 10542 7082
rect 10486 7028 10542 7030
rect 10590 7082 10646 7084
rect 10590 7030 10592 7082
rect 10592 7030 10644 7082
rect 10644 7030 10646 7082
rect 10590 7028 10646 7030
rect 11676 9660 11732 9716
rect 10892 6972 10948 7028
rect 11676 6972 11732 7028
rect 11116 6860 11172 6916
rect 10780 6748 10836 6804
rect 10332 6578 10388 6580
rect 10332 6526 10334 6578
rect 10334 6526 10386 6578
rect 10386 6526 10388 6578
rect 10332 6524 10388 6526
rect 10382 5514 10438 5516
rect 10382 5462 10384 5514
rect 10384 5462 10436 5514
rect 10436 5462 10438 5514
rect 10382 5460 10438 5462
rect 10486 5514 10542 5516
rect 10486 5462 10488 5514
rect 10488 5462 10540 5514
rect 10540 5462 10542 5514
rect 10486 5460 10542 5462
rect 10590 5514 10646 5516
rect 10590 5462 10592 5514
rect 10592 5462 10644 5514
rect 10644 5462 10646 5514
rect 10590 5460 10646 5462
rect 10220 4508 10276 4564
rect 11004 6412 11060 6468
rect 11004 5180 11060 5236
rect 10220 4172 10276 4228
rect 10108 3612 10164 3668
rect 10382 3946 10438 3948
rect 10382 3894 10384 3946
rect 10384 3894 10436 3946
rect 10436 3894 10438 3946
rect 10382 3892 10438 3894
rect 10486 3946 10542 3948
rect 10486 3894 10488 3946
rect 10488 3894 10540 3946
rect 10540 3894 10542 3946
rect 10486 3892 10542 3894
rect 10590 3946 10646 3948
rect 10590 3894 10592 3946
rect 10592 3894 10644 3946
rect 10644 3894 10646 3946
rect 10590 3892 10646 3894
rect 10220 3554 10276 3556
rect 10220 3502 10222 3554
rect 10222 3502 10274 3554
rect 10274 3502 10276 3554
rect 10220 3500 10276 3502
rect 10382 2378 10438 2380
rect 10382 2326 10384 2378
rect 10384 2326 10436 2378
rect 10436 2326 10438 2378
rect 10382 2324 10438 2326
rect 10486 2378 10542 2380
rect 10486 2326 10488 2378
rect 10488 2326 10540 2378
rect 10540 2326 10542 2378
rect 10486 2324 10542 2326
rect 10590 2378 10646 2380
rect 10590 2326 10592 2378
rect 10592 2326 10644 2378
rect 10644 2326 10646 2378
rect 10590 2324 10646 2326
rect 11452 4508 11508 4564
rect 11788 6748 11844 6804
rect 11788 5234 11844 5236
rect 11788 5182 11790 5234
rect 11790 5182 11842 5234
rect 11842 5182 11844 5234
rect 11788 5180 11844 5182
rect 12440 9434 12496 9436
rect 12440 9382 12442 9434
rect 12442 9382 12494 9434
rect 12494 9382 12496 9434
rect 12440 9380 12496 9382
rect 12544 9434 12600 9436
rect 12544 9382 12546 9434
rect 12546 9382 12598 9434
rect 12598 9382 12600 9434
rect 12544 9380 12600 9382
rect 12648 9434 12704 9436
rect 12648 9382 12650 9434
rect 12650 9382 12702 9434
rect 12702 9382 12704 9434
rect 12648 9380 12704 9382
rect 12796 8204 12852 8260
rect 12440 7866 12496 7868
rect 12440 7814 12442 7866
rect 12442 7814 12494 7866
rect 12494 7814 12496 7866
rect 12440 7812 12496 7814
rect 12544 7866 12600 7868
rect 12544 7814 12546 7866
rect 12546 7814 12598 7866
rect 12598 7814 12600 7866
rect 12544 7812 12600 7814
rect 12648 7866 12704 7868
rect 12648 7814 12650 7866
rect 12650 7814 12702 7866
rect 12702 7814 12704 7866
rect 12648 7812 12704 7814
rect 12236 7644 12292 7700
rect 13132 7644 13188 7700
rect 12124 6748 12180 6804
rect 12012 4284 12068 4340
rect 11788 3554 11844 3556
rect 11788 3502 11790 3554
rect 11790 3502 11842 3554
rect 11842 3502 11844 3554
rect 11788 3500 11844 3502
rect 11788 3276 11844 3332
rect 12012 3276 12068 3332
rect 12440 6298 12496 6300
rect 12440 6246 12442 6298
rect 12442 6246 12494 6298
rect 12494 6246 12496 6298
rect 12440 6244 12496 6246
rect 12544 6298 12600 6300
rect 12544 6246 12546 6298
rect 12546 6246 12598 6298
rect 12598 6246 12600 6298
rect 12544 6244 12600 6246
rect 12648 6298 12704 6300
rect 12648 6246 12650 6298
rect 12650 6246 12702 6298
rect 12702 6246 12704 6298
rect 12648 6244 12704 6246
rect 12796 5068 12852 5124
rect 12440 4730 12496 4732
rect 12440 4678 12442 4730
rect 12442 4678 12494 4730
rect 12494 4678 12496 4730
rect 12440 4676 12496 4678
rect 12544 4730 12600 4732
rect 12544 4678 12546 4730
rect 12546 4678 12598 4730
rect 12598 4678 12600 4730
rect 12544 4676 12600 4678
rect 12648 4730 12704 4732
rect 12648 4678 12650 4730
rect 12650 4678 12702 4730
rect 12702 4678 12704 4730
rect 12648 4676 12704 4678
rect 12684 4338 12740 4340
rect 12684 4286 12686 4338
rect 12686 4286 12738 4338
rect 12738 4286 12740 4338
rect 12684 4284 12740 4286
rect 12440 3162 12496 3164
rect 12440 3110 12442 3162
rect 12442 3110 12494 3162
rect 12494 3110 12496 3162
rect 12440 3108 12496 3110
rect 12544 3162 12600 3164
rect 12544 3110 12546 3162
rect 12546 3110 12598 3162
rect 12598 3110 12600 3162
rect 12544 3108 12600 3110
rect 12648 3162 12704 3164
rect 12648 3110 12650 3162
rect 12650 3110 12702 3162
rect 12702 3110 12704 3162
rect 12648 3108 12704 3110
rect 12440 1594 12496 1596
rect 12440 1542 12442 1594
rect 12442 1542 12494 1594
rect 12494 1542 12496 1594
rect 12440 1540 12496 1542
rect 12544 1594 12600 1596
rect 12544 1542 12546 1594
rect 12546 1542 12598 1594
rect 12598 1542 12600 1594
rect 12544 1540 12600 1542
rect 12648 1594 12704 1596
rect 12648 1542 12650 1594
rect 12650 1542 12702 1594
rect 12702 1542 12704 1594
rect 12648 1540 12704 1542
rect 13244 6636 13300 6692
rect 13468 5068 13524 5124
rect 13916 9100 13972 9156
rect 14498 10218 14554 10220
rect 14498 10166 14500 10218
rect 14500 10166 14552 10218
rect 14552 10166 14554 10218
rect 14498 10164 14554 10166
rect 14602 10218 14658 10220
rect 14602 10166 14604 10218
rect 14604 10166 14656 10218
rect 14656 10166 14658 10218
rect 14602 10164 14658 10166
rect 14706 10218 14762 10220
rect 14706 10166 14708 10218
rect 14708 10166 14760 10218
rect 14760 10166 14762 10218
rect 14706 10164 14762 10166
rect 14924 9884 14980 9940
rect 14924 9100 14980 9156
rect 14476 9042 14532 9044
rect 14476 8990 14478 9042
rect 14478 8990 14530 9042
rect 14530 8990 14532 9042
rect 14476 8988 14532 8990
rect 14498 8650 14554 8652
rect 14498 8598 14500 8650
rect 14500 8598 14552 8650
rect 14552 8598 14554 8650
rect 14498 8596 14554 8598
rect 14602 8650 14658 8652
rect 14602 8598 14604 8650
rect 14604 8598 14656 8650
rect 14656 8598 14658 8650
rect 14602 8596 14658 8598
rect 14706 8650 14762 8652
rect 14706 8598 14708 8650
rect 14708 8598 14760 8650
rect 14760 8598 14762 8650
rect 14706 8596 14762 8598
rect 14588 8258 14644 8260
rect 14588 8206 14590 8258
rect 14590 8206 14642 8258
rect 14642 8206 14644 8258
rect 14588 8204 14644 8206
rect 14140 7698 14196 7700
rect 14140 7646 14142 7698
rect 14142 7646 14194 7698
rect 14194 7646 14196 7698
rect 14140 7644 14196 7646
rect 14498 7082 14554 7084
rect 14498 7030 14500 7082
rect 14500 7030 14552 7082
rect 14552 7030 14554 7082
rect 14498 7028 14554 7030
rect 14602 7082 14658 7084
rect 14602 7030 14604 7082
rect 14604 7030 14656 7082
rect 14656 7030 14658 7082
rect 14602 7028 14658 7030
rect 14706 7082 14762 7084
rect 14706 7030 14708 7082
rect 14708 7030 14760 7082
rect 14760 7030 14762 7082
rect 14706 7028 14762 7030
rect 14588 6690 14644 6692
rect 14588 6638 14590 6690
rect 14590 6638 14642 6690
rect 14642 6638 14644 6690
rect 14588 6636 14644 6638
rect 14028 6188 14084 6244
rect 13692 4508 13748 4564
rect 13692 4338 13748 4340
rect 13692 4286 13694 4338
rect 13694 4286 13746 4338
rect 13746 4286 13748 4338
rect 13692 4284 13748 4286
rect 13692 3500 13748 3556
rect 13916 2098 13972 2100
rect 13916 2046 13918 2098
rect 13918 2046 13970 2098
rect 13970 2046 13972 2098
rect 13916 2044 13972 2046
rect 14140 3276 14196 3332
rect 14498 5514 14554 5516
rect 14498 5462 14500 5514
rect 14500 5462 14552 5514
rect 14552 5462 14554 5514
rect 14498 5460 14554 5462
rect 14602 5514 14658 5516
rect 14602 5462 14604 5514
rect 14604 5462 14656 5514
rect 14656 5462 14658 5514
rect 14602 5460 14658 5462
rect 14706 5514 14762 5516
rect 14706 5462 14708 5514
rect 14708 5462 14760 5514
rect 14760 5462 14762 5514
rect 14706 5460 14762 5462
rect 14498 3946 14554 3948
rect 14498 3894 14500 3946
rect 14500 3894 14552 3946
rect 14552 3894 14554 3946
rect 14498 3892 14554 3894
rect 14602 3946 14658 3948
rect 14602 3894 14604 3946
rect 14604 3894 14656 3946
rect 14656 3894 14658 3946
rect 14602 3892 14658 3894
rect 14706 3946 14762 3948
rect 14706 3894 14708 3946
rect 14708 3894 14760 3946
rect 14760 3894 14762 3946
rect 14706 3892 14762 3894
rect 14588 3554 14644 3556
rect 14588 3502 14590 3554
rect 14590 3502 14642 3554
rect 14642 3502 14644 3554
rect 14588 3500 14644 3502
rect 14476 2658 14532 2660
rect 14476 2606 14478 2658
rect 14478 2606 14530 2658
rect 14530 2606 14532 2658
rect 14476 2604 14532 2606
rect 14498 2378 14554 2380
rect 14498 2326 14500 2378
rect 14500 2326 14552 2378
rect 14552 2326 14554 2378
rect 14498 2324 14554 2326
rect 14602 2378 14658 2380
rect 14602 2326 14604 2378
rect 14604 2326 14656 2378
rect 14656 2326 14658 2378
rect 14602 2324 14658 2326
rect 14706 2378 14762 2380
rect 14706 2326 14708 2378
rect 14708 2326 14760 2378
rect 14760 2326 14762 2378
rect 14706 2324 14762 2326
rect 15036 6188 15092 6244
rect 15036 5180 15092 5236
rect 15484 9938 15540 9940
rect 15484 9886 15486 9938
rect 15486 9886 15538 9938
rect 15538 9886 15540 9938
rect 15484 9884 15540 9886
rect 15484 9042 15540 9044
rect 15484 8990 15486 9042
rect 15486 8990 15538 9042
rect 15538 8990 15540 9042
rect 15484 8988 15540 8990
rect 16268 9660 16324 9716
rect 16556 9434 16612 9436
rect 16556 9382 16558 9434
rect 16558 9382 16610 9434
rect 16610 9382 16612 9434
rect 16556 9380 16612 9382
rect 16660 9434 16716 9436
rect 16660 9382 16662 9434
rect 16662 9382 16714 9434
rect 16714 9382 16716 9434
rect 16660 9380 16716 9382
rect 16764 9434 16820 9436
rect 16764 9382 16766 9434
rect 16766 9382 16818 9434
rect 16818 9382 16820 9434
rect 16764 9380 16820 9382
rect 16156 8428 16212 8484
rect 15596 8258 15652 8260
rect 15596 8206 15598 8258
rect 15598 8206 15650 8258
rect 15650 8206 15652 8258
rect 15596 8204 15652 8206
rect 15596 6690 15652 6692
rect 15596 6638 15598 6690
rect 15598 6638 15650 6690
rect 15650 6638 15652 6690
rect 15596 6636 15652 6638
rect 15596 5234 15652 5236
rect 15596 5182 15598 5234
rect 15598 5182 15650 5234
rect 15650 5182 15652 5234
rect 15596 5180 15652 5182
rect 15596 3554 15652 3556
rect 15596 3502 15598 3554
rect 15598 3502 15650 3554
rect 15650 3502 15652 3554
rect 15596 3500 15652 3502
rect 15372 2604 15428 2660
rect 15036 1986 15092 1988
rect 15036 1934 15038 1986
rect 15038 1934 15090 1986
rect 15090 1934 15092 1986
rect 15036 1932 15092 1934
rect 15820 2044 15876 2100
rect 15596 1932 15652 1988
rect 16556 7866 16612 7868
rect 16556 7814 16558 7866
rect 16558 7814 16610 7866
rect 16610 7814 16612 7866
rect 16556 7812 16612 7814
rect 16660 7866 16716 7868
rect 16660 7814 16662 7866
rect 16662 7814 16714 7866
rect 16714 7814 16716 7866
rect 16660 7812 16716 7814
rect 16764 7866 16820 7868
rect 16764 7814 16766 7866
rect 16766 7814 16818 7866
rect 16818 7814 16820 7866
rect 16764 7812 16820 7814
rect 16556 6298 16612 6300
rect 16556 6246 16558 6298
rect 16558 6246 16610 6298
rect 16610 6246 16612 6298
rect 16556 6244 16612 6246
rect 16660 6298 16716 6300
rect 16660 6246 16662 6298
rect 16662 6246 16714 6298
rect 16714 6246 16716 6298
rect 16660 6244 16716 6246
rect 16764 6298 16820 6300
rect 16764 6246 16766 6298
rect 16766 6246 16818 6298
rect 16818 6246 16820 6298
rect 16764 6244 16820 6246
rect 16556 4730 16612 4732
rect 16556 4678 16558 4730
rect 16558 4678 16610 4730
rect 16610 4678 16612 4730
rect 16556 4676 16612 4678
rect 16660 4730 16716 4732
rect 16660 4678 16662 4730
rect 16662 4678 16714 4730
rect 16714 4678 16716 4730
rect 16660 4676 16716 4678
rect 16764 4730 16820 4732
rect 16764 4678 16766 4730
rect 16766 4678 16818 4730
rect 16818 4678 16820 4730
rect 16764 4676 16820 4678
rect 16556 3162 16612 3164
rect 16556 3110 16558 3162
rect 16558 3110 16610 3162
rect 16610 3110 16612 3162
rect 16556 3108 16612 3110
rect 16660 3162 16716 3164
rect 16660 3110 16662 3162
rect 16662 3110 16714 3162
rect 16714 3110 16716 3162
rect 16660 3108 16716 3110
rect 16764 3162 16820 3164
rect 16764 3110 16766 3162
rect 16766 3110 16818 3162
rect 16818 3110 16820 3162
rect 16764 3108 16820 3110
rect 16556 1594 16612 1596
rect 16556 1542 16558 1594
rect 16558 1542 16610 1594
rect 16610 1542 16612 1594
rect 16556 1540 16612 1542
rect 16660 1594 16716 1596
rect 16660 1542 16662 1594
rect 16662 1542 16714 1594
rect 16714 1542 16716 1594
rect 16660 1540 16716 1542
rect 16764 1594 16820 1596
rect 16764 1542 16766 1594
rect 16766 1542 16818 1594
rect 16818 1542 16820 1594
rect 16764 1540 16820 1542
<< metal3 >>
rect 2140 10164 2150 10220
rect 2206 10164 2254 10220
rect 2310 10164 2358 10220
rect 2414 10164 2424 10220
rect 6256 10164 6266 10220
rect 6322 10164 6370 10220
rect 6426 10164 6474 10220
rect 6530 10164 6540 10220
rect 10372 10164 10382 10220
rect 10438 10164 10486 10220
rect 10542 10164 10590 10220
rect 10646 10164 10656 10220
rect 14488 10164 14498 10220
rect 14554 10164 14602 10220
rect 14658 10164 14706 10220
rect 14762 10164 14772 10220
rect 14914 9884 14924 9940
rect 14980 9884 15484 9940
rect 15540 9884 15550 9940
rect 1586 9772 1596 9828
rect 1652 9772 3388 9828
rect 3444 9772 4956 9828
rect 5012 9772 5022 9828
rect 11666 9660 11676 9716
rect 11732 9660 16268 9716
rect 16324 9660 16334 9716
rect 4198 9380 4208 9436
rect 4264 9380 4312 9436
rect 4368 9380 4416 9436
rect 4472 9380 4482 9436
rect 8314 9380 8324 9436
rect 8380 9380 8428 9436
rect 8484 9380 8532 9436
rect 8588 9380 8598 9436
rect 12430 9380 12440 9436
rect 12496 9380 12544 9436
rect 12600 9380 12648 9436
rect 12704 9380 12714 9436
rect 16546 9380 16556 9436
rect 16612 9380 16660 9436
rect 16716 9380 16764 9436
rect 16820 9380 16830 9436
rect 13906 9100 13916 9156
rect 13972 9100 14924 9156
rect 14980 9100 14990 9156
rect 14466 8988 14476 9044
rect 14532 8988 15484 9044
rect 15540 8988 15550 9044
rect 0 8932 800 8960
rect 16200 8932 17000 8960
rect 0 8876 5068 8932
rect 5124 8876 5292 8932
rect 5348 8876 5358 8932
rect 8372 8876 17000 8932
rect 0 8848 800 8876
rect 8372 8820 8428 8876
rect 16200 8848 17000 8876
rect 7634 8764 7644 8820
rect 7700 8764 8428 8820
rect 2818 8652 2828 8708
rect 2884 8652 4396 8708
rect 4452 8652 4462 8708
rect 2140 8596 2150 8652
rect 2206 8596 2254 8652
rect 2310 8596 2358 8652
rect 2414 8596 2424 8652
rect 6256 8596 6266 8652
rect 6322 8596 6370 8652
rect 6426 8596 6474 8652
rect 6530 8596 6540 8652
rect 10372 8596 10382 8652
rect 10438 8596 10486 8652
rect 10542 8596 10590 8652
rect 10646 8596 10656 8652
rect 14488 8596 14498 8652
rect 14554 8596 14602 8652
rect 14658 8596 14706 8652
rect 14762 8596 14772 8652
rect 10770 8428 10780 8484
rect 10836 8428 16156 8484
rect 16212 8428 16222 8484
rect 12786 8204 12796 8260
rect 12852 8204 14588 8260
rect 14644 8204 15596 8260
rect 15652 8204 15662 8260
rect 2706 8092 2716 8148
rect 2772 8092 6076 8148
rect 6132 8092 6142 8148
rect 3490 7980 3500 8036
rect 3556 7980 4508 8036
rect 4564 7980 4574 8036
rect 4198 7812 4208 7868
rect 4264 7812 4312 7868
rect 4368 7812 4416 7868
rect 4472 7812 4482 7868
rect 8314 7812 8324 7868
rect 8380 7812 8428 7868
rect 8484 7812 8532 7868
rect 8588 7812 8598 7868
rect 12430 7812 12440 7868
rect 12496 7812 12544 7868
rect 12600 7812 12648 7868
rect 12704 7812 12714 7868
rect 16546 7812 16556 7868
rect 16612 7812 16660 7868
rect 16716 7812 16764 7868
rect 16820 7812 16830 7868
rect 12226 7644 12236 7700
rect 12292 7644 13132 7700
rect 13188 7644 14140 7700
rect 14196 7644 14206 7700
rect 6066 7532 6076 7588
rect 6132 7532 7308 7588
rect 7364 7532 7374 7588
rect 5058 7420 5068 7476
rect 5124 7420 6300 7476
rect 6356 7420 7364 7476
rect 7308 7364 7364 7420
rect 2594 7308 2604 7364
rect 2660 7308 4060 7364
rect 4116 7308 4126 7364
rect 7298 7308 7308 7364
rect 7364 7308 7374 7364
rect 2140 7028 2150 7084
rect 2206 7028 2254 7084
rect 2310 7028 2358 7084
rect 2414 7028 2424 7084
rect 6256 7028 6266 7084
rect 6322 7028 6370 7084
rect 6426 7028 6474 7084
rect 6530 7028 6540 7084
rect 10372 7028 10382 7084
rect 10438 7028 10486 7084
rect 10542 7028 10590 7084
rect 10646 7028 10656 7084
rect 14488 7028 14498 7084
rect 14554 7028 14602 7084
rect 14658 7028 14706 7084
rect 14762 7028 14772 7084
rect 10882 6972 10892 7028
rect 10948 6972 11676 7028
rect 11732 6972 11742 7028
rect 8642 6860 8652 6916
rect 8708 6860 11116 6916
rect 11172 6860 11182 6916
rect 9538 6748 9548 6804
rect 9604 6748 10780 6804
rect 10836 6748 10846 6804
rect 11778 6748 11788 6804
rect 11844 6748 12124 6804
rect 12180 6748 12190 6804
rect 2594 6636 2604 6692
rect 2660 6636 3388 6692
rect 3444 6636 5404 6692
rect 5460 6636 5470 6692
rect 7970 6636 7980 6692
rect 8036 6636 8876 6692
rect 8932 6636 9884 6692
rect 9940 6636 9950 6692
rect 13234 6636 13244 6692
rect 13300 6636 14588 6692
rect 14644 6636 15596 6692
rect 15652 6636 15662 6692
rect 1922 6524 1932 6580
rect 1988 6524 3500 6580
rect 3556 6524 3566 6580
rect 8194 6524 8204 6580
rect 8260 6524 9324 6580
rect 9380 6524 10332 6580
rect 10388 6524 10398 6580
rect 9986 6412 9996 6468
rect 10052 6412 11004 6468
rect 11060 6412 11070 6468
rect 4198 6244 4208 6300
rect 4264 6244 4312 6300
rect 4368 6244 4416 6300
rect 4472 6244 4482 6300
rect 8314 6244 8324 6300
rect 8380 6244 8428 6300
rect 8484 6244 8532 6300
rect 8588 6244 8598 6300
rect 12430 6244 12440 6300
rect 12496 6244 12544 6300
rect 12600 6244 12648 6300
rect 12704 6244 12714 6300
rect 16546 6244 16556 6300
rect 16612 6244 16660 6300
rect 16716 6244 16764 6300
rect 16820 6244 16830 6300
rect 14018 6188 14028 6244
rect 14084 6188 15036 6244
rect 15092 6188 15102 6244
rect 3154 5852 3164 5908
rect 3220 5852 4172 5908
rect 4228 5852 4956 5908
rect 5012 5852 5022 5908
rect 2140 5460 2150 5516
rect 2206 5460 2254 5516
rect 2310 5460 2358 5516
rect 2414 5460 2424 5516
rect 6256 5460 6266 5516
rect 6322 5460 6370 5516
rect 6426 5460 6474 5516
rect 6530 5460 6540 5516
rect 10372 5460 10382 5516
rect 10438 5460 10486 5516
rect 10542 5460 10590 5516
rect 10646 5460 10656 5516
rect 14488 5460 14498 5516
rect 14554 5460 14602 5516
rect 14658 5460 14706 5516
rect 14762 5460 14772 5516
rect 10994 5180 11004 5236
rect 11060 5180 11788 5236
rect 11844 5180 11854 5236
rect 15026 5180 15036 5236
rect 15092 5180 15596 5236
rect 15652 5180 15662 5236
rect 3826 5068 3836 5124
rect 3892 5068 4508 5124
rect 4564 5068 6636 5124
rect 6692 5068 6702 5124
rect 12786 5068 12796 5124
rect 12852 5068 13468 5124
rect 13524 5068 13534 5124
rect 1026 4956 1036 5012
rect 1092 4956 2492 5012
rect 2548 4956 2558 5012
rect 7196 4844 8988 4900
rect 9044 4844 9054 4900
rect 7196 4788 7252 4844
rect 5954 4732 5964 4788
rect 6020 4732 7196 4788
rect 7252 4732 7262 4788
rect 4198 4676 4208 4732
rect 4264 4676 4312 4732
rect 4368 4676 4416 4732
rect 4472 4676 4482 4732
rect 8314 4676 8324 4732
rect 8380 4676 8428 4732
rect 8484 4676 8532 4732
rect 8588 4676 8598 4732
rect 12430 4676 12440 4732
rect 12496 4676 12544 4732
rect 12600 4676 12648 4732
rect 12704 4676 12714 4732
rect 16546 4676 16556 4732
rect 16612 4676 16660 4732
rect 16716 4676 16764 4732
rect 16820 4676 16830 4732
rect 7858 4508 7868 4564
rect 7924 4508 10220 4564
rect 10276 4508 10286 4564
rect 11442 4508 11452 4564
rect 11508 4508 13692 4564
rect 13748 4508 13758 4564
rect 1474 4396 1484 4452
rect 1540 4396 3612 4452
rect 3668 4396 3678 4452
rect 4610 4284 4620 4340
rect 4676 4284 5852 4340
rect 5908 4284 6860 4340
rect 6916 4284 6926 4340
rect 12002 4284 12012 4340
rect 12068 4284 12684 4340
rect 12740 4284 13692 4340
rect 13748 4284 13758 4340
rect 9090 4172 9100 4228
rect 9156 4172 10220 4228
rect 10276 4172 10286 4228
rect 6850 4060 6860 4116
rect 6916 4060 7532 4116
rect 7588 4060 8540 4116
rect 8596 4060 8606 4116
rect 2140 3892 2150 3948
rect 2206 3892 2254 3948
rect 2310 3892 2358 3948
rect 2414 3892 2424 3948
rect 6256 3892 6266 3948
rect 6322 3892 6370 3948
rect 6426 3892 6474 3948
rect 6530 3892 6540 3948
rect 10372 3892 10382 3948
rect 10438 3892 10486 3948
rect 10542 3892 10590 3948
rect 10646 3892 10656 3948
rect 14488 3892 14498 3948
rect 14554 3892 14602 3948
rect 14658 3892 14706 3948
rect 14762 3892 14772 3948
rect 578 3612 588 3668
rect 644 3612 2380 3668
rect 2436 3612 2446 3668
rect 6514 3612 6524 3668
rect 6580 3612 10108 3668
rect 10164 3612 10174 3668
rect 10210 3500 10220 3556
rect 10276 3500 11788 3556
rect 11844 3500 11854 3556
rect 13682 3500 13692 3556
rect 13748 3500 14588 3556
rect 14644 3500 15596 3556
rect 15652 3500 15662 3556
rect 3266 3388 3276 3444
rect 3332 3388 3724 3444
rect 3780 3388 4508 3444
rect 4564 3388 4574 3444
rect 11778 3276 11788 3332
rect 11844 3276 12012 3332
rect 12068 3276 14140 3332
rect 14196 3276 14206 3332
rect 4198 3108 4208 3164
rect 4264 3108 4312 3164
rect 4368 3108 4416 3164
rect 4472 3108 4482 3164
rect 8314 3108 8324 3164
rect 8380 3108 8428 3164
rect 8484 3108 8532 3164
rect 8588 3108 8598 3164
rect 12430 3108 12440 3164
rect 12496 3108 12544 3164
rect 12600 3108 12648 3164
rect 12704 3108 12714 3164
rect 16546 3108 16556 3164
rect 16612 3108 16660 3164
rect 16716 3108 16764 3164
rect 16820 3108 16830 3164
rect 0 2996 800 3024
rect 16200 2996 17000 3024
rect 0 2940 1596 2996
rect 1652 2940 2156 2996
rect 2212 2940 2222 2996
rect 12348 2940 17000 2996
rect 0 2912 800 2940
rect 7298 2716 7308 2772
rect 7364 2716 8540 2772
rect 8596 2716 8606 2772
rect 12348 2660 12404 2940
rect 16200 2912 17000 2940
rect 4498 2604 4508 2660
rect 4564 2604 12404 2660
rect 14466 2604 14476 2660
rect 14532 2604 15372 2660
rect 15428 2604 15438 2660
rect 2140 2324 2150 2380
rect 2206 2324 2254 2380
rect 2310 2324 2358 2380
rect 2414 2324 2424 2380
rect 6256 2324 6266 2380
rect 6322 2324 6370 2380
rect 6426 2324 6474 2380
rect 6530 2324 6540 2380
rect 10372 2324 10382 2380
rect 10438 2324 10486 2380
rect 10542 2324 10590 2380
rect 10646 2324 10656 2380
rect 14488 2324 14498 2380
rect 14554 2324 14602 2380
rect 14658 2324 14706 2380
rect 14762 2324 14772 2380
rect 13906 2044 13916 2100
rect 13972 2044 15820 2100
rect 15876 2044 15886 2100
rect 15026 1932 15036 1988
rect 15092 1932 15596 1988
rect 15652 1932 15662 1988
rect 5506 1820 5516 1876
rect 5572 1820 6748 1876
rect 6804 1820 7756 1876
rect 7812 1820 7822 1876
rect 4198 1540 4208 1596
rect 4264 1540 4312 1596
rect 4368 1540 4416 1596
rect 4472 1540 4482 1596
rect 8314 1540 8324 1596
rect 8380 1540 8428 1596
rect 8484 1540 8532 1596
rect 8588 1540 8598 1596
rect 12430 1540 12440 1596
rect 12496 1540 12544 1596
rect 12600 1540 12648 1596
rect 12704 1540 12714 1596
rect 16546 1540 16556 1596
rect 16612 1540 16660 1596
rect 16716 1540 16764 1596
rect 16820 1540 16830 1596
<< via3 >>
rect 2150 10164 2206 10220
rect 2254 10164 2310 10220
rect 2358 10164 2414 10220
rect 6266 10164 6322 10220
rect 6370 10164 6426 10220
rect 6474 10164 6530 10220
rect 10382 10164 10438 10220
rect 10486 10164 10542 10220
rect 10590 10164 10646 10220
rect 14498 10164 14554 10220
rect 14602 10164 14658 10220
rect 14706 10164 14762 10220
rect 4208 9380 4264 9436
rect 4312 9380 4368 9436
rect 4416 9380 4472 9436
rect 8324 9380 8380 9436
rect 8428 9380 8484 9436
rect 8532 9380 8588 9436
rect 12440 9380 12496 9436
rect 12544 9380 12600 9436
rect 12648 9380 12704 9436
rect 16556 9380 16612 9436
rect 16660 9380 16716 9436
rect 16764 9380 16820 9436
rect 2150 8596 2206 8652
rect 2254 8596 2310 8652
rect 2358 8596 2414 8652
rect 6266 8596 6322 8652
rect 6370 8596 6426 8652
rect 6474 8596 6530 8652
rect 10382 8596 10438 8652
rect 10486 8596 10542 8652
rect 10590 8596 10646 8652
rect 14498 8596 14554 8652
rect 14602 8596 14658 8652
rect 14706 8596 14762 8652
rect 4208 7812 4264 7868
rect 4312 7812 4368 7868
rect 4416 7812 4472 7868
rect 8324 7812 8380 7868
rect 8428 7812 8484 7868
rect 8532 7812 8588 7868
rect 12440 7812 12496 7868
rect 12544 7812 12600 7868
rect 12648 7812 12704 7868
rect 16556 7812 16612 7868
rect 16660 7812 16716 7868
rect 16764 7812 16820 7868
rect 2150 7028 2206 7084
rect 2254 7028 2310 7084
rect 2358 7028 2414 7084
rect 6266 7028 6322 7084
rect 6370 7028 6426 7084
rect 6474 7028 6530 7084
rect 10382 7028 10438 7084
rect 10486 7028 10542 7084
rect 10590 7028 10646 7084
rect 14498 7028 14554 7084
rect 14602 7028 14658 7084
rect 14706 7028 14762 7084
rect 4208 6244 4264 6300
rect 4312 6244 4368 6300
rect 4416 6244 4472 6300
rect 8324 6244 8380 6300
rect 8428 6244 8484 6300
rect 8532 6244 8588 6300
rect 12440 6244 12496 6300
rect 12544 6244 12600 6300
rect 12648 6244 12704 6300
rect 16556 6244 16612 6300
rect 16660 6244 16716 6300
rect 16764 6244 16820 6300
rect 2150 5460 2206 5516
rect 2254 5460 2310 5516
rect 2358 5460 2414 5516
rect 6266 5460 6322 5516
rect 6370 5460 6426 5516
rect 6474 5460 6530 5516
rect 10382 5460 10438 5516
rect 10486 5460 10542 5516
rect 10590 5460 10646 5516
rect 14498 5460 14554 5516
rect 14602 5460 14658 5516
rect 14706 5460 14762 5516
rect 4208 4676 4264 4732
rect 4312 4676 4368 4732
rect 4416 4676 4472 4732
rect 8324 4676 8380 4732
rect 8428 4676 8484 4732
rect 8532 4676 8588 4732
rect 12440 4676 12496 4732
rect 12544 4676 12600 4732
rect 12648 4676 12704 4732
rect 16556 4676 16612 4732
rect 16660 4676 16716 4732
rect 16764 4676 16820 4732
rect 2150 3892 2206 3948
rect 2254 3892 2310 3948
rect 2358 3892 2414 3948
rect 6266 3892 6322 3948
rect 6370 3892 6426 3948
rect 6474 3892 6530 3948
rect 10382 3892 10438 3948
rect 10486 3892 10542 3948
rect 10590 3892 10646 3948
rect 14498 3892 14554 3948
rect 14602 3892 14658 3948
rect 14706 3892 14762 3948
rect 4208 3108 4264 3164
rect 4312 3108 4368 3164
rect 4416 3108 4472 3164
rect 8324 3108 8380 3164
rect 8428 3108 8484 3164
rect 8532 3108 8588 3164
rect 12440 3108 12496 3164
rect 12544 3108 12600 3164
rect 12648 3108 12704 3164
rect 16556 3108 16612 3164
rect 16660 3108 16716 3164
rect 16764 3108 16820 3164
rect 2150 2324 2206 2380
rect 2254 2324 2310 2380
rect 2358 2324 2414 2380
rect 6266 2324 6322 2380
rect 6370 2324 6426 2380
rect 6474 2324 6530 2380
rect 10382 2324 10438 2380
rect 10486 2324 10542 2380
rect 10590 2324 10646 2380
rect 14498 2324 14554 2380
rect 14602 2324 14658 2380
rect 14706 2324 14762 2380
rect 4208 1540 4264 1596
rect 4312 1540 4368 1596
rect 4416 1540 4472 1596
rect 8324 1540 8380 1596
rect 8428 1540 8484 1596
rect 8532 1540 8588 1596
rect 12440 1540 12496 1596
rect 12544 1540 12600 1596
rect 12648 1540 12704 1596
rect 16556 1540 16612 1596
rect 16660 1540 16716 1596
rect 16764 1540 16820 1596
<< metal4 >>
rect 2122 10220 2442 10252
rect 2122 10164 2150 10220
rect 2206 10164 2254 10220
rect 2310 10164 2358 10220
rect 2414 10164 2442 10220
rect 2122 8652 2442 10164
rect 2122 8596 2150 8652
rect 2206 8596 2254 8652
rect 2310 8596 2358 8652
rect 2414 8596 2442 8652
rect 2122 7084 2442 8596
rect 2122 7028 2150 7084
rect 2206 7028 2254 7084
rect 2310 7028 2358 7084
rect 2414 7028 2442 7084
rect 2122 5516 2442 7028
rect 2122 5460 2150 5516
rect 2206 5460 2254 5516
rect 2310 5460 2358 5516
rect 2414 5460 2442 5516
rect 2122 3948 2442 5460
rect 2122 3892 2150 3948
rect 2206 3892 2254 3948
rect 2310 3892 2358 3948
rect 2414 3892 2442 3948
rect 2122 2380 2442 3892
rect 2122 2324 2150 2380
rect 2206 2324 2254 2380
rect 2310 2324 2358 2380
rect 2414 2324 2442 2380
rect 2122 1508 2442 2324
rect 4180 9436 4500 10252
rect 4180 9380 4208 9436
rect 4264 9380 4312 9436
rect 4368 9380 4416 9436
rect 4472 9380 4500 9436
rect 4180 7868 4500 9380
rect 4180 7812 4208 7868
rect 4264 7812 4312 7868
rect 4368 7812 4416 7868
rect 4472 7812 4500 7868
rect 4180 6300 4500 7812
rect 4180 6244 4208 6300
rect 4264 6244 4312 6300
rect 4368 6244 4416 6300
rect 4472 6244 4500 6300
rect 4180 4732 4500 6244
rect 4180 4676 4208 4732
rect 4264 4676 4312 4732
rect 4368 4676 4416 4732
rect 4472 4676 4500 4732
rect 4180 3164 4500 4676
rect 4180 3108 4208 3164
rect 4264 3108 4312 3164
rect 4368 3108 4416 3164
rect 4472 3108 4500 3164
rect 4180 1596 4500 3108
rect 4180 1540 4208 1596
rect 4264 1540 4312 1596
rect 4368 1540 4416 1596
rect 4472 1540 4500 1596
rect 4180 1508 4500 1540
rect 6238 10220 6558 10252
rect 6238 10164 6266 10220
rect 6322 10164 6370 10220
rect 6426 10164 6474 10220
rect 6530 10164 6558 10220
rect 6238 8652 6558 10164
rect 6238 8596 6266 8652
rect 6322 8596 6370 8652
rect 6426 8596 6474 8652
rect 6530 8596 6558 8652
rect 6238 7084 6558 8596
rect 6238 7028 6266 7084
rect 6322 7028 6370 7084
rect 6426 7028 6474 7084
rect 6530 7028 6558 7084
rect 6238 5516 6558 7028
rect 6238 5460 6266 5516
rect 6322 5460 6370 5516
rect 6426 5460 6474 5516
rect 6530 5460 6558 5516
rect 6238 3948 6558 5460
rect 6238 3892 6266 3948
rect 6322 3892 6370 3948
rect 6426 3892 6474 3948
rect 6530 3892 6558 3948
rect 6238 2380 6558 3892
rect 6238 2324 6266 2380
rect 6322 2324 6370 2380
rect 6426 2324 6474 2380
rect 6530 2324 6558 2380
rect 6238 1508 6558 2324
rect 8296 9436 8616 10252
rect 8296 9380 8324 9436
rect 8380 9380 8428 9436
rect 8484 9380 8532 9436
rect 8588 9380 8616 9436
rect 8296 7868 8616 9380
rect 8296 7812 8324 7868
rect 8380 7812 8428 7868
rect 8484 7812 8532 7868
rect 8588 7812 8616 7868
rect 8296 6300 8616 7812
rect 8296 6244 8324 6300
rect 8380 6244 8428 6300
rect 8484 6244 8532 6300
rect 8588 6244 8616 6300
rect 8296 4732 8616 6244
rect 8296 4676 8324 4732
rect 8380 4676 8428 4732
rect 8484 4676 8532 4732
rect 8588 4676 8616 4732
rect 8296 3164 8616 4676
rect 8296 3108 8324 3164
rect 8380 3108 8428 3164
rect 8484 3108 8532 3164
rect 8588 3108 8616 3164
rect 8296 1596 8616 3108
rect 8296 1540 8324 1596
rect 8380 1540 8428 1596
rect 8484 1540 8532 1596
rect 8588 1540 8616 1596
rect 8296 1508 8616 1540
rect 10354 10220 10674 10252
rect 10354 10164 10382 10220
rect 10438 10164 10486 10220
rect 10542 10164 10590 10220
rect 10646 10164 10674 10220
rect 10354 8652 10674 10164
rect 10354 8596 10382 8652
rect 10438 8596 10486 8652
rect 10542 8596 10590 8652
rect 10646 8596 10674 8652
rect 10354 7084 10674 8596
rect 10354 7028 10382 7084
rect 10438 7028 10486 7084
rect 10542 7028 10590 7084
rect 10646 7028 10674 7084
rect 10354 5516 10674 7028
rect 10354 5460 10382 5516
rect 10438 5460 10486 5516
rect 10542 5460 10590 5516
rect 10646 5460 10674 5516
rect 10354 3948 10674 5460
rect 10354 3892 10382 3948
rect 10438 3892 10486 3948
rect 10542 3892 10590 3948
rect 10646 3892 10674 3948
rect 10354 2380 10674 3892
rect 10354 2324 10382 2380
rect 10438 2324 10486 2380
rect 10542 2324 10590 2380
rect 10646 2324 10674 2380
rect 10354 1508 10674 2324
rect 12412 9436 12732 10252
rect 12412 9380 12440 9436
rect 12496 9380 12544 9436
rect 12600 9380 12648 9436
rect 12704 9380 12732 9436
rect 12412 7868 12732 9380
rect 12412 7812 12440 7868
rect 12496 7812 12544 7868
rect 12600 7812 12648 7868
rect 12704 7812 12732 7868
rect 12412 6300 12732 7812
rect 12412 6244 12440 6300
rect 12496 6244 12544 6300
rect 12600 6244 12648 6300
rect 12704 6244 12732 6300
rect 12412 4732 12732 6244
rect 12412 4676 12440 4732
rect 12496 4676 12544 4732
rect 12600 4676 12648 4732
rect 12704 4676 12732 4732
rect 12412 3164 12732 4676
rect 12412 3108 12440 3164
rect 12496 3108 12544 3164
rect 12600 3108 12648 3164
rect 12704 3108 12732 3164
rect 12412 1596 12732 3108
rect 12412 1540 12440 1596
rect 12496 1540 12544 1596
rect 12600 1540 12648 1596
rect 12704 1540 12732 1596
rect 12412 1508 12732 1540
rect 14470 10220 14790 10252
rect 14470 10164 14498 10220
rect 14554 10164 14602 10220
rect 14658 10164 14706 10220
rect 14762 10164 14790 10220
rect 14470 8652 14790 10164
rect 14470 8596 14498 8652
rect 14554 8596 14602 8652
rect 14658 8596 14706 8652
rect 14762 8596 14790 8652
rect 14470 7084 14790 8596
rect 14470 7028 14498 7084
rect 14554 7028 14602 7084
rect 14658 7028 14706 7084
rect 14762 7028 14790 7084
rect 14470 5516 14790 7028
rect 14470 5460 14498 5516
rect 14554 5460 14602 5516
rect 14658 5460 14706 5516
rect 14762 5460 14790 5516
rect 14470 3948 14790 5460
rect 14470 3892 14498 3948
rect 14554 3892 14602 3948
rect 14658 3892 14706 3948
rect 14762 3892 14790 3948
rect 14470 2380 14790 3892
rect 14470 2324 14498 2380
rect 14554 2324 14602 2380
rect 14658 2324 14706 2380
rect 14762 2324 14790 2380
rect 14470 1508 14790 2324
rect 16528 9436 16848 10252
rect 16528 9380 16556 9436
rect 16612 9380 16660 9436
rect 16716 9380 16764 9436
rect 16820 9380 16848 9436
rect 16528 7868 16848 9380
rect 16528 7812 16556 7868
rect 16612 7812 16660 7868
rect 16716 7812 16764 7868
rect 16820 7812 16848 7868
rect 16528 6300 16848 7812
rect 16528 6244 16556 6300
rect 16612 6244 16660 6300
rect 16716 6244 16764 6300
rect 16820 6244 16848 6300
rect 16528 4732 16848 6244
rect 16528 4676 16556 4732
rect 16612 4676 16660 4732
rect 16716 4676 16764 4732
rect 16820 4676 16848 4732
rect 16528 3164 16848 4676
rect 16528 3108 16556 3164
rect 16612 3108 16660 3164
rect 16716 3108 16764 3164
rect 16820 3108 16848 3164
rect 16528 1596 16848 3108
rect 16528 1540 16556 1596
rect 16612 1540 16660 1596
rect 16716 1540 16764 1596
rect 16820 1540 16848 1596
rect 16528 1508 16848 1540
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_BUF\[0\]_I OpenLane/pdks/gf180mcuC/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1666464484
transform 1 0 11536 0 1 1568
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_BUF\[1\]_I
timestamp 1666464484
transform 1 0 11760 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_BUF\[2\]_I
timestamp 1666464484
transform 1 0 11312 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_BUF\[3\]_I
timestamp 1666464484
transform 1 0 11760 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_BUF\[4\]_I
timestamp 1666464484
transform 1 0 7840 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_BUF\[5\]_I
timestamp 1666464484
transform 1 0 14112 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_BUF\[6\]_I
timestamp 1666464484
transform 1 0 11760 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_BUF\[7\]_I
timestamp 1666464484
transform 1 0 13664 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_BUF\[8\]_I
timestamp 1666464484
transform 1 0 14112 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_BUF\[9\]_I
timestamp 1666464484
transform 1 0 15568 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_BUF\[10\]_I
timestamp 1666464484
transform 1 0 15568 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_BUF\[11\]_I
timestamp 1666464484
transform 1 0 15568 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_BUF\[12\]_I
timestamp 1666464484
transform 1 0 15568 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_BUF\[13\]_I
timestamp 1666464484
transform 1 0 15456 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_BUF\[14\]_I
timestamp 1666464484
transform 1 0 15456 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_BUF\[15\]_I
timestamp 1666464484
transform 1 0 16016 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_BUF\[16\]_I
timestamp 1666464484
transform -1 0 15680 0 1 1568
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_BUF\[17\]_I
timestamp 1666464484
transform -1 0 11984 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_BUF\[18\]_I
timestamp 1666464484
transform 1 0 1568 0 -1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_BUF\[19\]_I
timestamp 1666464484
transform -1 0 5152 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_BUF\[20\]_I
timestamp 1666464484
transform 1 0 672 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_BUF\[21\]_I
timestamp 1666464484
transform -1 0 896 0 1 1568
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_BUF\[22\]_I
timestamp 1666464484
transform 1 0 5040 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_BUF\[23\]_I
timestamp 1666464484
transform 1 0 4480 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_BUF\[24\]_I
timestamp 1666464484
transform 1 0 5376 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_BUF\[25\]_I
timestamp 1666464484
transform 1 0 4592 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_BUF\[26\]_I
timestamp 1666464484
transform 1 0 4928 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_BUF\[27\]_I
timestamp 1666464484
transform 1 0 4480 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_BUF\[28\]_I
timestamp 1666464484
transform 1 0 4480 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_BUF\[29\]_I
timestamp 1666464484
transform 1 0 6832 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_BUF\[30\]_I
timestamp 1666464484
transform 1 0 7280 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_BUF\[31\]_I
timestamp 1666464484
transform 1 0 7728 0 1 1568
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_BUF\[32\]_I
timestamp 1666464484
transform 1 0 8960 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_BUF\[33\]_I
timestamp 1666464484
transform 1 0 4480 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_BUF\[34\]_I
timestamp 1666464484
transform 1 0 8512 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_BUF\[35\]_I
timestamp 1666464484
transform 1 0 8512 0 -1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_BUF\[36\]_I
timestamp 1666464484
transform 1 0 9856 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_BUF\[37\]_I
timestamp 1666464484
transform 1 0 10304 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_8  BUF\[0\] OpenLane/pdks/gf180mcuC/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1666464484
transform -1 0 11312 0 1 1568
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_8  BUF\[1\]
timestamp 1666464484
transform -1 0 10976 0 1 3136
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_8  BUF\[2\]
timestamp 1666464484
transform -1 0 11312 0 1 4704
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_8  BUF\[3\]
timestamp 1666464484
transform -1 0 11760 0 -1 6272
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_8  BUF\[4\]
timestamp 1666464484
transform -1 0 7840 0 1 3136
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_8  BUF\[5\]
timestamp 1666464484
transform -1 0 12656 0 -1 3136
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_8  BUF\[6\]
timestamp 1666464484
transform 1 0 11984 0 -1 6272
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_8  BUF\[7\]
timestamp 1666464484
transform -1 0 13440 0 -1 4704
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_8  BUF\[8\]
timestamp 1666464484
transform -1 0 13888 0 -1 7840
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_8  BUF\[9\]
timestamp 1666464484
transform -1 0 15344 0 1 7840
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_8  BUF\[10\]
timestamp 1666464484
transform -1 0 15344 0 1 6272
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_8  BUF\[11\]
timestamp 1666464484
transform -1 0 15344 0 1 3136
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_8  BUF\[12\]
timestamp 1666464484
transform -1 0 15344 0 1 4704
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_8  BUF\[13\]
timestamp 1666464484
transform -1 0 15232 0 -1 9408
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_8  BUF\[14\]
timestamp 1666464484
transform -1 0 15232 0 1 9408
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_8  BUF\[15\]
timestamp 1666464484
transform -1 0 15792 0 -1 3136
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_8  BUF\[16\]
timestamp 1666464484
transform -1 0 15232 0 1 1568
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_8  BUF\[17\]
timestamp 1666464484
transform -1 0 12096 0 -1 9408
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_8  BUF\[18\]
timestamp 1666464484
transform 1 0 2016 0 -1 3136
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_8  BUF\[19\]
timestamp 1666464484
transform 1 0 5152 0 -1 9408
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_8  BUF\[20\]
timestamp 1666464484
transform 1 0 1120 0 1 3136
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_8  BUF\[21\]
timestamp 1666464484
transform 1 0 1120 0 1 1568
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_8  BUF\[22\]
timestamp 1666464484
transform -1 0 4032 0 1 9408
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_8  BUF\[23\]
timestamp 1666464484
transform -1 0 4032 0 1 7840
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_8  BUF\[24\]
timestamp 1666464484
transform -1 0 4032 0 1 6272
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_8  BUF\[25\]
timestamp 1666464484
transform -1 0 4592 0 -1 9408
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_8  BUF\[26\]
timestamp 1666464484
transform -1 0 4928 0 -1 6272
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_8  BUF\[27\]
timestamp 1666464484
transform -1 0 3472 0 -1 4704
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_8  BUF\[28\]
timestamp 1666464484
transform -1 0 3920 0 -1 7840
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_8  BUF\[29\]
timestamp 1666464484
transform -1 0 6608 0 -1 4704
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_8  BUF\[30\]
timestamp 1666464484
transform -1 0 7056 0 -1 7840
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_8  BUF\[31\]
timestamp 1666464484
transform -1 0 7504 0 1 1568
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_8  BUF\[32\]
timestamp 1666464484
transform -1 0 7952 0 1 4704
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_8  BUF\[33\]
timestamp 1666464484
transform -1 0 4032 0 1 4704
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_8  BUF\[34\]
timestamp 1666464484
transform -1 0 8064 0 -1 6272
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_8  BUF\[35\]
timestamp 1666464484
transform -1 0 8064 0 -1 3136
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_8  BUF\[36\]
timestamp 1666464484
transform -1 0 9632 0 1 7840
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_8  BUF\[37\]
timestamp 1666464484
transform -1 0 10080 0 1 6272
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_2 OpenLane/pdks/gf180mcuC/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1666464484
transform 1 0 448 0 1 1568
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_6
timestamp 1666464484
transform 1 0 896 0 1 1568
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_34 OpenLane/pdks/gf180mcuC/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1666464484
transform 1 0 4032 0 1 1568
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_37
timestamp 1666464484
transform 1 0 4368 0 1 1568
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_65
timestamp 1666464484
transform 1 0 7504 0 1 1568
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_69
timestamp 1666464484
transform 1 0 7952 0 1 1568
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_72
timestamp 1666464484
transform 1 0 8288 0 1 1568
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_99
timestamp 1666464484
transform 1 0 11312 0 1 1568
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_103
timestamp 1666464484
transform 1 0 11760 0 1 1568
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_107
timestamp 1666464484
transform 1 0 12208 0 1 1568
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_134
timestamp 1666464484
transform 1 0 15232 0 1 1568
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_138
timestamp 1666464484
transform 1 0 15680 0 1 1568
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_142
timestamp 1666464484
transform 1 0 16128 0 1 1568
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_144
timestamp 1666464484
transform 1 0 16352 0 1 1568
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_1_2 OpenLane/pdks/gf180mcuC/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1666464484
transform 1 0 448 0 -1 3136
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_1_10
timestamp 1666464484
transform 1 0 1344 0 -1 3136
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_1_14
timestamp 1666464484
transform 1 0 1792 0 -1 3136
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_1_42
timestamp 1666464484
transform 1 0 4928 0 -1 3136
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_1_70
timestamp 1666464484
transform 1 0 8064 0 -1 3136
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_1_73
timestamp 1666464484
transform 1 0 8400 0 -1 3136
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_1_76
timestamp 1666464484
transform 1 0 8736 0 -1 3136
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_1_84
timestamp 1666464484
transform 1 0 9632 0 -1 3136
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_1_111
timestamp 1666464484
transform 1 0 12656 0 -1 3136
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_1_139
timestamp 1666464484
transform 1 0 15792 0 -1 3136
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_1_141
timestamp 1666464484
transform 1 0 16016 0 -1 3136
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_1_144
timestamp 1666464484
transform 1 0 16352 0 -1 3136
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_2_2
timestamp 1666464484
transform 1 0 448 0 1 3136
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_2_6
timestamp 1666464484
transform 1 0 896 0 1 3136
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_2_34
timestamp 1666464484
transform 1 0 4032 0 1 3136
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_2_37
timestamp 1666464484
transform 1 0 4368 0 1 3136
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_2_40
timestamp 1666464484
transform 1 0 4704 0 1 3136
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_2_68
timestamp 1666464484
transform 1 0 7840 0 1 3136
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_2_96
timestamp 1666464484
transform 1 0 10976 0 1 3136
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_2_98
timestamp 1666464484
transform 1 0 11200 0 1 3136
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_2_101
timestamp 1666464484
transform 1 0 11536 0 1 3136
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_2_105
timestamp 1666464484
transform 1 0 11984 0 1 3136
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_2_108
timestamp 1666464484
transform 1 0 12320 0 1 3136
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_2_135
timestamp 1666464484
transform 1 0 15344 0 1 3136
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_2_139
timestamp 1666464484
transform 1 0 15792 0 1 3136
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_2_143
timestamp 1666464484
transform 1 0 16240 0 1 3136
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_3_2
timestamp 1666464484
transform 1 0 448 0 -1 4704
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_3_29
timestamp 1666464484
transform 1 0 3472 0 -1 4704
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_3_57
timestamp 1666464484
transform 1 0 6608 0 -1 4704
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_3_61 OpenLane/pdks/gf180mcuC/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1666464484
transform 1 0 7056 0 -1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_3_65
timestamp 1666464484
transform 1 0 7504 0 -1 4704
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_3_67
timestamp 1666464484
transform 1 0 7728 0 -1 4704
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_3_70
timestamp 1666464484
transform 1 0 8064 0 -1 4704
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_3_73
timestamp 1666464484
transform 1 0 8400 0 -1 4704
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_3_76
timestamp 1666464484
transform 1 0 8736 0 -1 4704
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_3_80
timestamp 1666464484
transform 1 0 9184 0 -1 4704
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_3_88
timestamp 1666464484
transform 1 0 10080 0 -1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_3_118
timestamp 1666464484
transform 1 0 13440 0 -1 4704
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_3_122
timestamp 1666464484
transform 1 0 13888 0 -1 4704
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_3_126 OpenLane/pdks/gf180mcuC/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1666464484
transform 1 0 14336 0 -1 4704
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_3_144
timestamp 1666464484
transform 1 0 16352 0 -1 4704
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_4_2
timestamp 1666464484
transform 1 0 448 0 1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_4_6
timestamp 1666464484
transform 1 0 896 0 1 4704
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_4_34
timestamp 1666464484
transform 1 0 4032 0 1 4704
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_4_37
timestamp 1666464484
transform 1 0 4368 0 1 4704
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_4_40
timestamp 1666464484
transform 1 0 4704 0 1 4704
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_4_42
timestamp 1666464484
transform 1 0 4928 0 1 4704
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_4_69
timestamp 1666464484
transform 1 0 7952 0 1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_4_99
timestamp 1666464484
transform 1 0 11312 0 1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_4_105
timestamp 1666464484
transform 1 0 11984 0 1 4704
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_4_108
timestamp 1666464484
transform 1 0 12320 0 1 4704
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_4_135
timestamp 1666464484
transform 1 0 15344 0 1 4704
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_4_139
timestamp 1666464484
transform 1 0 15792 0 1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_4_143
timestamp 1666464484
transform 1 0 16240 0 1 4704
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_5_2
timestamp 1666464484
transform 1 0 448 0 -1 6272
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_5_10
timestamp 1666464484
transform 1 0 1344 0 -1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_5_14
timestamp 1666464484
transform 1 0 1792 0 -1 6272
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_5_42
timestamp 1666464484
transform 1 0 4928 0 -1 6272
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_5_70
timestamp 1666464484
transform 1 0 8064 0 -1 6272
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_5_73
timestamp 1666464484
transform 1 0 8400 0 -1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_5_103
timestamp 1666464484
transform 1 0 11760 0 -1 6272
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_5_131
timestamp 1666464484
transform 1 0 14896 0 -1 6272
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_5_139
timestamp 1666464484
transform 1 0 15792 0 -1 6272
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_5_141
timestamp 1666464484
transform 1 0 16016 0 -1 6272
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_5_144
timestamp 1666464484
transform 1 0 16352 0 -1 6272
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_6_2
timestamp 1666464484
transform 1 0 448 0 1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_6_6
timestamp 1666464484
transform 1 0 896 0 1 6272
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_6_34
timestamp 1666464484
transform 1 0 4032 0 1 6272
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_6_37
timestamp 1666464484
transform 1 0 4368 0 1 6272
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_6_40
timestamp 1666464484
transform 1 0 4704 0 1 6272
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_6_44
timestamp 1666464484
transform 1 0 5152 0 1 6272
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_6_48
timestamp 1666464484
transform 1 0 5600 0 1 6272
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_6_56
timestamp 1666464484
transform 1 0 6496 0 1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_6_60
timestamp 1666464484
transform 1 0 6944 0 1 6272
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_6_88
timestamp 1666464484
transform 1 0 10080 0 1 6272
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_6_92
timestamp 1666464484
transform 1 0 10528 0 1 6272
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_6_100
timestamp 1666464484
transform 1 0 11424 0 1 6272
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_6_102
timestamp 1666464484
transform 1 0 11648 0 1 6272
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_6_105
timestamp 1666464484
transform 1 0 11984 0 1 6272
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_6_108
timestamp 1666464484
transform 1 0 12320 0 1 6272
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_6_135
timestamp 1666464484
transform 1 0 15344 0 1 6272
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_6_139
timestamp 1666464484
transform 1 0 15792 0 1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_6_143
timestamp 1666464484
transform 1 0 16240 0 1 6272
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_7_2
timestamp 1666464484
transform 1 0 448 0 -1 7840
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_7_6
timestamp 1666464484
transform 1 0 896 0 -1 7840
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_7_33
timestamp 1666464484
transform 1 0 3920 0 -1 7840
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_7_61
timestamp 1666464484
transform 1 0 7056 0 -1 7840
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_7_65
timestamp 1666464484
transform 1 0 7504 0 -1 7840
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_7_69
timestamp 1666464484
transform 1 0 7952 0 -1 7840
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_7_73
timestamp 1666464484
transform 1 0 8400 0 -1 7840
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_7_89
timestamp 1666464484
transform 1 0 10192 0 -1 7840
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_7_93
timestamp 1666464484
transform 1 0 10640 0 -1 7840
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_7_95
timestamp 1666464484
transform 1 0 10864 0 -1 7840
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_7_122
timestamp 1666464484
transform 1 0 13888 0 -1 7840
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_7_126
timestamp 1666464484
transform 1 0 14336 0 -1 7840
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_7_144
timestamp 1666464484
transform 1 0 16352 0 -1 7840
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_8_2
timestamp 1666464484
transform 1 0 448 0 1 7840
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_8_6
timestamp 1666464484
transform 1 0 896 0 1 7840
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_8_34
timestamp 1666464484
transform 1 0 4032 0 1 7840
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_8_37
timestamp 1666464484
transform 1 0 4368 0 1 7840
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_8_40
timestamp 1666464484
transform 1 0 4704 0 1 7840
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_8_44
timestamp 1666464484
transform 1 0 5152 0 1 7840
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_8_52
timestamp 1666464484
transform 1 0 6048 0 1 7840
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_8_56
timestamp 1666464484
transform 1 0 6496 0 1 7840
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_8_84
timestamp 1666464484
transform 1 0 9632 0 1 7840
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_8_88
timestamp 1666464484
transform 1 0 10080 0 1 7840
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_8_96
timestamp 1666464484
transform 1 0 10976 0 1 7840
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_8_100
timestamp 1666464484
transform 1 0 11424 0 1 7840
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_8_102
timestamp 1666464484
transform 1 0 11648 0 1 7840
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_8_105
timestamp 1666464484
transform 1 0 11984 0 1 7840
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_8_108
timestamp 1666464484
transform 1 0 12320 0 1 7840
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_8_135
timestamp 1666464484
transform 1 0 15344 0 1 7840
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_8_139
timestamp 1666464484
transform 1 0 15792 0 1 7840
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_8_143
timestamp 1666464484
transform 1 0 16240 0 1 7840
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_9_2
timestamp 1666464484
transform 1 0 448 0 -1 9408
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_9_10
timestamp 1666464484
transform 1 0 1344 0 -1 9408
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_9_12
timestamp 1666464484
transform 1 0 1568 0 -1 9408
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_9_39
timestamp 1666464484
transform 1 0 4592 0 -1 9408
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_9_43
timestamp 1666464484
transform 1 0 5040 0 -1 9408
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_9_70
timestamp 1666464484
transform 1 0 8064 0 -1 9408
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_9_73
timestamp 1666464484
transform 1 0 8400 0 -1 9408
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_9_77
timestamp 1666464484
transform 1 0 8848 0 -1 9408
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_9_79
timestamp 1666464484
transform 1 0 9072 0 -1 9408
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_9_106
timestamp 1666464484
transform 1 0 12096 0 -1 9408
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_9_134
timestamp 1666464484
transform 1 0 15232 0 -1 9408
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_9_138
timestamp 1666464484
transform 1 0 15680 0 -1 9408
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_9_144
timestamp 1666464484
transform 1 0 16352 0 -1 9408
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_10_2
timestamp 1666464484
transform 1 0 448 0 1 9408
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_10_6
timestamp 1666464484
transform 1 0 896 0 1 9408
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_10_34
timestamp 1666464484
transform 1 0 4032 0 1 9408
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_10_37
timestamp 1666464484
transform 1 0 4368 0 1 9408
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_10_41
timestamp 1666464484
transform 1 0 4816 0 1 9408
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_10_45
timestamp 1666464484
transform 1 0 5264 0 1 9408
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_10_61
timestamp 1666464484
transform 1 0 7056 0 1 9408
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_10_69
timestamp 1666464484
transform 1 0 7952 0 1 9408
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_10_72 OpenLane/pdks/gf180mcuC/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1666464484
transform 1 0 8288 0 1 9408
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_10_104
timestamp 1666464484
transform 1 0 11872 0 1 9408
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_10_107
timestamp 1666464484
transform 1 0 12208 0 1 9408
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_10_134
timestamp 1666464484
transform 1 0 15232 0 1 9408
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_10_138
timestamp 1666464484
transform 1 0 15680 0 1 9408
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_10_142
timestamp 1666464484
transform 1 0 16128 0 1 9408
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_10_144
timestamp 1666464484
transform 1 0 16352 0 1 9408
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_0 OpenLane/pdks/gf180mcuC/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1666464484
transform 1 0 224 0 1 1568
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_1
timestamp 1666464484
transform -1 0 16688 0 1 1568
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_2
timestamp 1666464484
transform 1 0 224 0 -1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_3
timestamp 1666464484
transform -1 0 16688 0 -1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_4
timestamp 1666464484
transform 1 0 224 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_5
timestamp 1666464484
transform -1 0 16688 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_6
timestamp 1666464484
transform 1 0 224 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_7
timestamp 1666464484
transform -1 0 16688 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_8
timestamp 1666464484
transform 1 0 224 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_9
timestamp 1666464484
transform -1 0 16688 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_10
timestamp 1666464484
transform 1 0 224 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_11
timestamp 1666464484
transform -1 0 16688 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_12
timestamp 1666464484
transform 1 0 224 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_13
timestamp 1666464484
transform -1 0 16688 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_14
timestamp 1666464484
transform 1 0 224 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_15
timestamp 1666464484
transform -1 0 16688 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_16
timestamp 1666464484
transform 1 0 224 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_17
timestamp 1666464484
transform -1 0 16688 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_18
timestamp 1666464484
transform 1 0 224 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_19
timestamp 1666464484
transform -1 0 16688 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_20
timestamp 1666464484
transform 1 0 224 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_21
timestamp 1666464484
transform -1 0 16688 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_22 OpenLane/pdks/gf180mcuC/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1666464484
transform 1 0 4144 0 1 1568
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_23
timestamp 1666464484
transform 1 0 8064 0 1 1568
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_24
timestamp 1666464484
transform 1 0 11984 0 1 1568
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_25
timestamp 1666464484
transform 1 0 15904 0 1 1568
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_26
timestamp 1666464484
transform 1 0 8176 0 -1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_27
timestamp 1666464484
transform 1 0 16128 0 -1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_28
timestamp 1666464484
transform 1 0 4144 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_29
timestamp 1666464484
transform 1 0 12096 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_30
timestamp 1666464484
transform 1 0 8176 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_31
timestamp 1666464484
transform 1 0 16128 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_32
timestamp 1666464484
transform 1 0 4144 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_33
timestamp 1666464484
transform 1 0 12096 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_34
timestamp 1666464484
transform 1 0 8176 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_35
timestamp 1666464484
transform 1 0 16128 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_36
timestamp 1666464484
transform 1 0 4144 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_37
timestamp 1666464484
transform 1 0 12096 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_38
timestamp 1666464484
transform 1 0 8176 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_39
timestamp 1666464484
transform 1 0 16128 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_40
timestamp 1666464484
transform 1 0 4144 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_41
timestamp 1666464484
transform 1 0 12096 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_42
timestamp 1666464484
transform 1 0 8176 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_43
timestamp 1666464484
transform 1 0 16128 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_44
timestamp 1666464484
transform 1 0 4144 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_45
timestamp 1666464484
transform 1 0 8064 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_46
timestamp 1666464484
transform 1 0 11984 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_47
timestamp 1666464484
transform 1 0 15904 0 1 9408
box -86 -86 310 870
<< labels >>
flabel metal4 s 2122 1508 2442 10252 0 FreeSans 1280 90 0 0 VDD
port 0 nsew power bidirectional
flabel metal4 s 6238 1508 6558 10252 0 FreeSans 1280 90 0 0 VDD
port 0 nsew power bidirectional
flabel metal4 s 10354 1508 10674 10252 0 FreeSans 1280 90 0 0 VDD
port 0 nsew power bidirectional
flabel metal4 s 14470 1508 14790 10252 0 FreeSans 1280 90 0 0 VDD
port 0 nsew power bidirectional
flabel metal4 s 4180 1508 4500 10252 0 FreeSans 1280 90 0 0 VSS
port 1 nsew ground bidirectional
flabel metal4 s 8296 1508 8616 10252 0 FreeSans 1280 90 0 0 VSS
port 1 nsew ground bidirectional
flabel metal4 s 12412 1508 12732 10252 0 FreeSans 1280 90 0 0 VSS
port 1 nsew ground bidirectional
flabel metal4 s 16528 1508 16848 10252 0 FreeSans 1280 90 0 0 VSS
port 1 nsew ground bidirectional
flabel metal2 s 560 0 672 800 0 FreeSans 448 90 0 0 mgmt_gpio_in[0]
port 2 nsew signal input
flabel metal2 s 5040 0 5152 800 0 FreeSans 448 90 0 0 mgmt_gpio_in[10]
port 3 nsew signal input
flabel metal2 s 5488 0 5600 800 0 FreeSans 448 90 0 0 mgmt_gpio_in[11]
port 4 nsew signal input
flabel metal2 s 5936 0 6048 800 0 FreeSans 448 90 0 0 mgmt_gpio_in[12]
port 5 nsew signal input
flabel metal2 s 6384 0 6496 800 0 FreeSans 448 90 0 0 mgmt_gpio_in[13]
port 6 nsew signal input
flabel metal2 s 6832 0 6944 800 0 FreeSans 448 90 0 0 mgmt_gpio_in[14]
port 7 nsew signal input
flabel metal2 s 7280 0 7392 800 0 FreeSans 448 90 0 0 mgmt_gpio_in[15]
port 8 nsew signal input
flabel metal2 s 7728 0 7840 800 0 FreeSans 448 90 0 0 mgmt_gpio_in[16]
port 9 nsew signal input
flabel metal2 s 8176 0 8288 800 0 FreeSans 448 90 0 0 mgmt_gpio_in[17]
port 10 nsew signal input
flabel metal2 s 1008 0 1120 800 0 FreeSans 448 90 0 0 mgmt_gpio_in[1]
port 11 nsew signal input
flabel metal2 s 1456 0 1568 800 0 FreeSans 448 90 0 0 mgmt_gpio_in[2]
port 12 nsew signal input
flabel metal2 s 1904 0 2016 800 0 FreeSans 448 90 0 0 mgmt_gpio_in[3]
port 13 nsew signal input
flabel metal2 s 2352 0 2464 800 0 FreeSans 448 90 0 0 mgmt_gpio_in[4]
port 14 nsew signal input
flabel metal2 s 2800 0 2912 800 0 FreeSans 448 90 0 0 mgmt_gpio_in[5]
port 15 nsew signal input
flabel metal2 s 3248 0 3360 800 0 FreeSans 448 90 0 0 mgmt_gpio_in[6]
port 16 nsew signal input
flabel metal2 s 3696 0 3808 800 0 FreeSans 448 90 0 0 mgmt_gpio_in[7]
port 17 nsew signal input
flabel metal2 s 4144 0 4256 800 0 FreeSans 448 90 0 0 mgmt_gpio_in[8]
port 18 nsew signal input
flabel metal2 s 4592 0 4704 800 0 FreeSans 448 90 0 0 mgmt_gpio_in[9]
port 19 nsew signal input
flabel metal2 s 560 11200 672 12000 0 FreeSans 448 90 0 0 mgmt_gpio_in_buf[0]
port 20 nsew signal tristate
flabel metal2 s 5040 11200 5152 12000 0 FreeSans 448 90 0 0 mgmt_gpio_in_buf[10]
port 21 nsew signal tristate
flabel metal2 s 5488 11200 5600 12000 0 FreeSans 448 90 0 0 mgmt_gpio_in_buf[11]
port 22 nsew signal tristate
flabel metal2 s 5936 11200 6048 12000 0 FreeSans 448 90 0 0 mgmt_gpio_in_buf[12]
port 23 nsew signal tristate
flabel metal2 s 6384 11200 6496 12000 0 FreeSans 448 90 0 0 mgmt_gpio_in_buf[13]
port 24 nsew signal tristate
flabel metal2 s 6832 11200 6944 12000 0 FreeSans 448 90 0 0 mgmt_gpio_in_buf[14]
port 25 nsew signal tristate
flabel metal2 s 7280 11200 7392 12000 0 FreeSans 448 90 0 0 mgmt_gpio_in_buf[15]
port 26 nsew signal tristate
flabel metal2 s 7728 11200 7840 12000 0 FreeSans 448 90 0 0 mgmt_gpio_in_buf[16]
port 27 nsew signal tristate
flabel metal2 s 8176 11200 8288 12000 0 FreeSans 448 90 0 0 mgmt_gpio_in_buf[17]
port 28 nsew signal tristate
flabel metal2 s 1008 11200 1120 12000 0 FreeSans 448 90 0 0 mgmt_gpio_in_buf[1]
port 29 nsew signal tristate
flabel metal2 s 1456 11200 1568 12000 0 FreeSans 448 90 0 0 mgmt_gpio_in_buf[2]
port 30 nsew signal tristate
flabel metal2 s 1904 11200 2016 12000 0 FreeSans 448 90 0 0 mgmt_gpio_in_buf[3]
port 31 nsew signal tristate
flabel metal2 s 2352 11200 2464 12000 0 FreeSans 448 90 0 0 mgmt_gpio_in_buf[4]
port 32 nsew signal tristate
flabel metal2 s 2800 11200 2912 12000 0 FreeSans 448 90 0 0 mgmt_gpio_in_buf[5]
port 33 nsew signal tristate
flabel metal2 s 3248 11200 3360 12000 0 FreeSans 448 90 0 0 mgmt_gpio_in_buf[6]
port 34 nsew signal tristate
flabel metal2 s 3696 11200 3808 12000 0 FreeSans 448 90 0 0 mgmt_gpio_in_buf[7]
port 35 nsew signal tristate
flabel metal2 s 4144 11200 4256 12000 0 FreeSans 448 90 0 0 mgmt_gpio_in_buf[8]
port 36 nsew signal tristate
flabel metal2 s 4592 11200 4704 12000 0 FreeSans 448 90 0 0 mgmt_gpio_in_buf[9]
port 37 nsew signal tristate
flabel metal3 s 0 2912 800 3024 0 FreeSans 448 0 0 0 mgmt_gpio_oeb[0]
port 38 nsew signal input
flabel metal3 s 0 8848 800 8960 0 FreeSans 448 0 0 0 mgmt_gpio_oeb[1]
port 39 nsew signal input
flabel metal3 s 16200 2912 17000 3024 0 FreeSans 448 0 0 0 mgmt_gpio_oeb_buf[0]
port 40 nsew signal tristate
flabel metal3 s 16200 8848 17000 8960 0 FreeSans 448 0 0 0 mgmt_gpio_oeb_buf[1]
port 41 nsew signal tristate
flabel metal2 s 8624 11200 8736 12000 0 FreeSans 448 90 0 0 mgmt_gpio_out[0]
port 42 nsew signal input
flabel metal2 s 13104 11200 13216 12000 0 FreeSans 448 90 0 0 mgmt_gpio_out[10]
port 43 nsew signal input
flabel metal2 s 13552 11200 13664 12000 0 FreeSans 448 90 0 0 mgmt_gpio_out[11]
port 44 nsew signal input
flabel metal2 s 14000 11200 14112 12000 0 FreeSans 448 90 0 0 mgmt_gpio_out[12]
port 45 nsew signal input
flabel metal2 s 14448 11200 14560 12000 0 FreeSans 448 90 0 0 mgmt_gpio_out[13]
port 46 nsew signal input
flabel metal2 s 14896 11200 15008 12000 0 FreeSans 448 90 0 0 mgmt_gpio_out[14]
port 47 nsew signal input
flabel metal2 s 15344 11200 15456 12000 0 FreeSans 448 90 0 0 mgmt_gpio_out[15]
port 48 nsew signal input
flabel metal2 s 15792 11200 15904 12000 0 FreeSans 448 90 0 0 mgmt_gpio_out[16]
port 49 nsew signal input
flabel metal2 s 16240 11200 16352 12000 0 FreeSans 448 90 0 0 mgmt_gpio_out[17]
port 50 nsew signal input
flabel metal2 s 9072 11200 9184 12000 0 FreeSans 448 90 0 0 mgmt_gpio_out[1]
port 51 nsew signal input
flabel metal2 s 9520 11200 9632 12000 0 FreeSans 448 90 0 0 mgmt_gpio_out[2]
port 52 nsew signal input
flabel metal2 s 9968 11200 10080 12000 0 FreeSans 448 90 0 0 mgmt_gpio_out[3]
port 53 nsew signal input
flabel metal2 s 10416 11200 10528 12000 0 FreeSans 448 90 0 0 mgmt_gpio_out[4]
port 54 nsew signal input
flabel metal2 s 10864 11200 10976 12000 0 FreeSans 448 90 0 0 mgmt_gpio_out[5]
port 55 nsew signal input
flabel metal2 s 11312 11200 11424 12000 0 FreeSans 448 90 0 0 mgmt_gpio_out[6]
port 56 nsew signal input
flabel metal2 s 11760 11200 11872 12000 0 FreeSans 448 90 0 0 mgmt_gpio_out[7]
port 57 nsew signal input
flabel metal2 s 12208 11200 12320 12000 0 FreeSans 448 90 0 0 mgmt_gpio_out[8]
port 58 nsew signal input
flabel metal2 s 12656 11200 12768 12000 0 FreeSans 448 90 0 0 mgmt_gpio_out[9]
port 59 nsew signal input
flabel metal2 s 8624 0 8736 800 0 FreeSans 448 90 0 0 mgmt_gpio_out_buf[0]
port 60 nsew signal tristate
flabel metal2 s 13104 0 13216 800 0 FreeSans 448 90 0 0 mgmt_gpio_out_buf[10]
port 61 nsew signal tristate
flabel metal2 s 13552 0 13664 800 0 FreeSans 448 90 0 0 mgmt_gpio_out_buf[11]
port 62 nsew signal tristate
flabel metal2 s 14000 0 14112 800 0 FreeSans 448 90 0 0 mgmt_gpio_out_buf[12]
port 63 nsew signal tristate
flabel metal2 s 14448 0 14560 800 0 FreeSans 448 90 0 0 mgmt_gpio_out_buf[13]
port 64 nsew signal tristate
flabel metal2 s 14896 0 15008 800 0 FreeSans 448 90 0 0 mgmt_gpio_out_buf[14]
port 65 nsew signal tristate
flabel metal2 s 15344 0 15456 800 0 FreeSans 448 90 0 0 mgmt_gpio_out_buf[15]
port 66 nsew signal tristate
flabel metal2 s 15792 0 15904 800 0 FreeSans 448 90 0 0 mgmt_gpio_out_buf[16]
port 67 nsew signal tristate
flabel metal2 s 16240 0 16352 800 0 FreeSans 448 90 0 0 mgmt_gpio_out_buf[17]
port 68 nsew signal tristate
flabel metal2 s 9072 0 9184 800 0 FreeSans 448 90 0 0 mgmt_gpio_out_buf[1]
port 69 nsew signal tristate
flabel metal2 s 9520 0 9632 800 0 FreeSans 448 90 0 0 mgmt_gpio_out_buf[2]
port 70 nsew signal tristate
flabel metal2 s 9968 0 10080 800 0 FreeSans 448 90 0 0 mgmt_gpio_out_buf[3]
port 71 nsew signal tristate
flabel metal2 s 10416 0 10528 800 0 FreeSans 448 90 0 0 mgmt_gpio_out_buf[4]
port 72 nsew signal tristate
flabel metal2 s 10864 0 10976 800 0 FreeSans 448 90 0 0 mgmt_gpio_out_buf[5]
port 73 nsew signal tristate
flabel metal2 s 11312 0 11424 800 0 FreeSans 448 90 0 0 mgmt_gpio_out_buf[6]
port 74 nsew signal tristate
flabel metal2 s 11760 0 11872 800 0 FreeSans 448 90 0 0 mgmt_gpio_out_buf[7]
port 75 nsew signal tristate
flabel metal2 s 12208 0 12320 800 0 FreeSans 448 90 0 0 mgmt_gpio_out_buf[8]
port 76 nsew signal tristate
flabel metal2 s 12656 0 12768 800 0 FreeSans 448 90 0 0 mgmt_gpio_out_buf[9]
port 77 nsew signal tristate
rlabel metal1 8456 10192 8456 10192 0 VDD
rlabel via1 8536 9408 8536 9408 0 VSS
rlabel metal2 672 3416 672 3416 0 mgmt_gpio_in[0]
rlabel metal3 5712 7448 5712 7448 0 mgmt_gpio_in[10]
rlabel metal2 6776 1904 6776 1904 0 mgmt_gpio_in[11]
rlabel metal2 7224 4928 7224 4928 0 mgmt_gpio_in[12]
rlabel metal3 5600 5096 5600 5096 0 mgmt_gpio_in[13]
rlabel metal2 6888 2422 6888 2422 0 mgmt_gpio_in[14]
rlabel metal2 7336 1750 7336 1750 0 mgmt_gpio_in[15]
rlabel metal2 7784 1190 7784 1190 0 mgmt_gpio_in[16]
rlabel metal2 8232 3654 8232 3654 0 mgmt_gpio_in[17]
rlabel metal2 1064 1960 1064 1960 0 mgmt_gpio_in[1]
rlabel metal2 1512 2366 1512 2366 0 mgmt_gpio_in[2]
rlabel metal2 3528 7392 3528 7392 0 mgmt_gpio_in[3]
rlabel metal3 3024 6664 3024 6664 0 mgmt_gpio_in[4]
rlabel metal2 4536 9016 4536 9016 0 mgmt_gpio_in[5]
rlabel metal3 3696 5880 3696 5880 0 mgmt_gpio_in[6]
rlabel metal3 4144 3416 4144 3416 0 mgmt_gpio_in[7]
rlabel metal2 4312 6440 4312 6440 0 mgmt_gpio_in[8]
rlabel metal3 5264 4312 5264 4312 0 mgmt_gpio_in[9]
rlabel metal3 1512 3640 1512 3640 0 mgmt_gpio_in_buf[0]
rlabel metal2 5152 9800 5152 9800 0 mgmt_gpio_in_buf[10]
rlabel metal2 5544 6650 5544 6650 0 mgmt_gpio_in_buf[11]
rlabel metal2 5992 8218 5992 8218 0 mgmt_gpio_in_buf[12]
rlabel metal3 4424 8120 4424 8120 0 mgmt_gpio_in_buf[13]
rlabel metal2 6664 7084 6664 7084 0 mgmt_gpio_in_buf[14]
rlabel metal3 6720 7560 6720 7560 0 mgmt_gpio_in_buf[15]
rlabel metal2 7784 9786 7784 9786 0 mgmt_gpio_in_buf[16]
rlabel metal2 8232 9002 8232 9002 0 mgmt_gpio_in_buf[17]
rlabel metal3 1792 4984 1792 4984 0 mgmt_gpio_in_buf[1]
rlabel metal2 1512 10570 1512 10570 0 mgmt_gpio_in_buf[2]
rlabel metal2 1960 9786 1960 9786 0 mgmt_gpio_in_buf[3]
rlabel metal2 2464 10360 2464 10360 0 mgmt_gpio_in_buf[4]
rlabel metal2 2856 10066 2856 10066 0 mgmt_gpio_in_buf[5]
rlabel metal2 3192 10024 3192 10024 0 mgmt_gpio_in_buf[6]
rlabel metal3 2576 4424 2576 4424 0 mgmt_gpio_in_buf[7]
rlabel metal3 3360 7336 3360 7336 0 mgmt_gpio_in_buf[8]
rlabel metal2 4704 9800 4704 9800 0 mgmt_gpio_in_buf[9]
rlabel metal3 1190 2968 1190 2968 0 mgmt_gpio_oeb[0]
rlabel metal3 2926 8904 2926 8904 0 mgmt_gpio_oeb[1]
rlabel metal3 12376 2800 12376 2800 0 mgmt_gpio_oeb_buf[0]
rlabel metal2 7672 8848 7672 8848 0 mgmt_gpio_oeb_buf[1]
rlabel metal2 11144 4424 11144 4424 0 mgmt_gpio_out[0]
rlabel metal3 13944 6664 13944 6664 0 mgmt_gpio_out[10]
rlabel metal3 14168 3528 14168 3528 0 mgmt_gpio_out[11]
rlabel metal2 15064 5656 15064 5656 0 mgmt_gpio_out[12]
rlabel metal2 14448 9016 14448 9016 0 mgmt_gpio_out[13]
rlabel metal2 14952 10514 14952 10514 0 mgmt_gpio_out[14]
rlabel metal2 16072 3696 16072 3696 0 mgmt_gpio_out[15]
rlabel metal2 15680 2072 15680 2072 0 mgmt_gpio_out[16]
rlabel metal2 11704 9352 11704 9352 0 mgmt_gpio_out[17]
rlabel metal2 10248 3864 10248 3864 0 mgmt_gpio_out[1]
rlabel metal2 10808 5936 10808 5936 0 mgmt_gpio_out[2]
rlabel metal2 11032 6160 11032 6160 0 mgmt_gpio_out[3]
rlabel metal2 7672 4032 7672 4032 0 mgmt_gpio_out[4]
rlabel metal2 12040 3024 12040 3024 0 mgmt_gpio_out[5]
rlabel metal2 12152 6328 12152 6328 0 mgmt_gpio_out[6]
rlabel metal3 12376 4312 12376 4312 0 mgmt_gpio_out[7]
rlabel metal2 13160 7560 13160 7560 0 mgmt_gpio_out[8]
rlabel metal3 13720 8232 13720 8232 0 mgmt_gpio_out[9]
rlabel metal2 8680 1414 8680 1414 0 mgmt_gpio_out_buf[0]
rlabel metal2 13160 3766 13160 3766 0 mgmt_gpio_out_buf[10]
rlabel metal2 13608 2198 13608 2198 0 mgmt_gpio_out_buf[11]
rlabel metal2 14056 2982 14056 2982 0 mgmt_gpio_out_buf[12]
rlabel metal2 14504 1246 14504 1246 0 mgmt_gpio_out_buf[13]
rlabel metal3 14448 9128 14448 9128 0 mgmt_gpio_out_buf[14]
rlabel metal2 15400 1694 15400 1694 0 mgmt_gpio_out_buf[15]
rlabel metal2 15848 1414 15848 1414 0 mgmt_gpio_out_buf[16]
rlabel metal2 16296 4578 16296 4578 0 mgmt_gpio_out_buf[17]
rlabel metal2 9128 2198 9128 2198 0 mgmt_gpio_out_buf[1]
rlabel metal2 9576 2982 9576 2982 0 mgmt_gpio_out_buf[2]
rlabel metal2 10024 3262 10024 3262 0 mgmt_gpio_out_buf[3]
rlabel metal2 10472 1302 10472 1302 0 mgmt_gpio_out_buf[4]
rlabel metal2 10920 1694 10920 1694 0 mgmt_gpio_out_buf[5]
rlabel metal2 11368 1806 11368 1806 0 mgmt_gpio_out_buf[6]
rlabel metal2 11816 1862 11816 1862 0 mgmt_gpio_out_buf[7]
rlabel metal2 12264 4046 12264 4046 0 mgmt_gpio_out_buf[8]
rlabel metal2 12712 1078 12712 1078 0 mgmt_gpio_out_buf[9]
<< properties >>
string FIXED_BBOX 0 0 17000 12000
<< end >>
