magic
tech gf180mcuC
magscale 1 5
timestamp 1668625752
<< obsm1 >>
rect 672 1538 46975 73401
<< metal2 >>
rect 2184 74600 2240 75000
rect 2800 74600 2856 75000
rect 3416 74600 3472 75000
rect 4032 74600 4088 75000
rect 4648 74600 4704 75000
rect 5264 74600 5320 75000
rect 5880 74600 5936 75000
rect 6496 74600 6552 75000
rect 7112 74600 7168 75000
rect 7728 74600 7784 75000
rect 8344 74600 8400 75000
rect 8960 74600 9016 75000
rect 9576 74600 9632 75000
rect 10192 74600 10248 75000
rect 10808 74600 10864 75000
rect 11424 74600 11480 75000
rect 12040 74600 12096 75000
rect 12656 74600 12712 75000
rect 13272 74600 13328 75000
rect 13888 74600 13944 75000
rect 14504 74600 14560 75000
rect 15120 74600 15176 75000
rect 15736 74600 15792 75000
rect 16352 74600 16408 75000
rect 16968 74600 17024 75000
rect 17584 74600 17640 75000
rect 18200 74600 18256 75000
rect 18816 74600 18872 75000
rect 19432 74600 19488 75000
rect 20048 74600 20104 75000
rect 20664 74600 20720 75000
rect 21280 74600 21336 75000
rect 21896 74600 21952 75000
rect 22512 74600 22568 75000
rect 23128 74600 23184 75000
rect 23744 74600 23800 75000
rect 24360 74600 24416 75000
rect 24976 74600 25032 75000
rect 25592 74600 25648 75000
rect 26208 74600 26264 75000
rect 26824 74600 26880 75000
rect 27440 74600 27496 75000
rect 28056 74600 28112 75000
rect 28672 74600 28728 75000
rect 29288 74600 29344 75000
rect 29904 74600 29960 75000
rect 30520 74600 30576 75000
rect 31136 74600 31192 75000
rect 31752 74600 31808 75000
rect 32368 74600 32424 75000
rect 32984 74600 33040 75000
rect 33600 74600 33656 75000
rect 34216 74600 34272 75000
rect 34832 74600 34888 75000
rect 35448 74600 35504 75000
rect 36064 74600 36120 75000
rect 36680 74600 36736 75000
rect 37296 74600 37352 75000
rect 37912 74600 37968 75000
rect 38528 74600 38584 75000
rect 39144 74600 39200 75000
rect 39760 74600 39816 75000
rect 40376 74600 40432 75000
rect 40992 74600 41048 75000
rect 41608 74600 41664 75000
rect 42224 74600 42280 75000
rect 42840 74600 42896 75000
rect 43456 74600 43512 75000
rect 44072 74600 44128 75000
rect 44688 74600 44744 75000
rect 1008 0 1064 400
rect 1512 0 1568 400
rect 2016 0 2072 400
rect 2520 0 2576 400
rect 3024 0 3080 400
rect 3528 0 3584 400
rect 4032 0 4088 400
rect 4536 0 4592 400
rect 5040 0 5096 400
rect 5544 0 5600 400
rect 6048 0 6104 400
rect 6552 0 6608 400
rect 7056 0 7112 400
rect 7560 0 7616 400
rect 8064 0 8120 400
rect 8568 0 8624 400
rect 9072 0 9128 400
rect 9576 0 9632 400
rect 10080 0 10136 400
rect 10584 0 10640 400
rect 11088 0 11144 400
rect 11592 0 11648 400
rect 12096 0 12152 400
rect 12600 0 12656 400
rect 13104 0 13160 400
rect 13608 0 13664 400
rect 14112 0 14168 400
rect 14616 0 14672 400
rect 15120 0 15176 400
rect 15624 0 15680 400
rect 16128 0 16184 400
rect 16632 0 16688 400
rect 17136 0 17192 400
rect 17640 0 17696 400
rect 18144 0 18200 400
rect 18648 0 18704 400
rect 19152 0 19208 400
rect 19656 0 19712 400
rect 20160 0 20216 400
rect 20664 0 20720 400
rect 21168 0 21224 400
rect 21672 0 21728 400
rect 22176 0 22232 400
rect 22680 0 22736 400
rect 23184 0 23240 400
rect 23688 0 23744 400
rect 24192 0 24248 400
rect 24696 0 24752 400
rect 25200 0 25256 400
rect 25704 0 25760 400
rect 26208 0 26264 400
rect 26712 0 26768 400
rect 27216 0 27272 400
rect 27720 0 27776 400
rect 28224 0 28280 400
rect 28728 0 28784 400
rect 29232 0 29288 400
rect 29736 0 29792 400
rect 30240 0 30296 400
rect 30744 0 30800 400
rect 31248 0 31304 400
rect 31752 0 31808 400
rect 32256 0 32312 400
rect 32760 0 32816 400
rect 33264 0 33320 400
rect 33768 0 33824 400
rect 34272 0 34328 400
rect 34776 0 34832 400
rect 35280 0 35336 400
rect 35784 0 35840 400
rect 36288 0 36344 400
rect 36792 0 36848 400
rect 37296 0 37352 400
rect 37800 0 37856 400
rect 38304 0 38360 400
rect 38808 0 38864 400
rect 39312 0 39368 400
rect 39816 0 39872 400
rect 40320 0 40376 400
rect 40824 0 40880 400
rect 41328 0 41384 400
rect 41832 0 41888 400
rect 42336 0 42392 400
rect 42840 0 42896 400
rect 43344 0 43400 400
rect 43848 0 43904 400
rect 44352 0 44408 400
rect 44856 0 44912 400
rect 45360 0 45416 400
rect 45864 0 45920 400
<< obsm2 >>
rect 742 74570 2154 74975
rect 2270 74570 2770 74975
rect 2886 74570 3386 74975
rect 3502 74570 4002 74975
rect 4118 74570 4618 74975
rect 4734 74570 5234 74975
rect 5350 74570 5850 74975
rect 5966 74570 6466 74975
rect 6582 74570 7082 74975
rect 7198 74570 7698 74975
rect 7814 74570 8314 74975
rect 8430 74570 8930 74975
rect 9046 74570 9546 74975
rect 9662 74570 10162 74975
rect 10278 74570 10778 74975
rect 10894 74570 11394 74975
rect 11510 74570 12010 74975
rect 12126 74570 12626 74975
rect 12742 74570 13242 74975
rect 13358 74570 13858 74975
rect 13974 74570 14474 74975
rect 14590 74570 15090 74975
rect 15206 74570 15706 74975
rect 15822 74570 16322 74975
rect 16438 74570 16938 74975
rect 17054 74570 17554 74975
rect 17670 74570 18170 74975
rect 18286 74570 18786 74975
rect 18902 74570 19402 74975
rect 19518 74570 20018 74975
rect 20134 74570 20634 74975
rect 20750 74570 21250 74975
rect 21366 74570 21866 74975
rect 21982 74570 22482 74975
rect 22598 74570 23098 74975
rect 23214 74570 23714 74975
rect 23830 74570 24330 74975
rect 24446 74570 24946 74975
rect 25062 74570 25562 74975
rect 25678 74570 26178 74975
rect 26294 74570 26794 74975
rect 26910 74570 27410 74975
rect 27526 74570 28026 74975
rect 28142 74570 28642 74975
rect 28758 74570 29258 74975
rect 29374 74570 29874 74975
rect 29990 74570 30490 74975
rect 30606 74570 31106 74975
rect 31222 74570 31722 74975
rect 31838 74570 32338 74975
rect 32454 74570 32954 74975
rect 33070 74570 33570 74975
rect 33686 74570 34186 74975
rect 34302 74570 34802 74975
rect 34918 74570 35418 74975
rect 35534 74570 36034 74975
rect 36150 74570 36650 74975
rect 36766 74570 37266 74975
rect 37382 74570 37882 74975
rect 37998 74570 38498 74975
rect 38614 74570 39114 74975
rect 39230 74570 39730 74975
rect 39846 74570 40346 74975
rect 40462 74570 40962 74975
rect 41078 74570 41578 74975
rect 41694 74570 42194 74975
rect 42310 74570 42810 74975
rect 42926 74570 43426 74975
rect 43542 74570 44042 74975
rect 44158 74570 44658 74975
rect 44774 74570 46970 74975
rect 742 430 46970 74570
rect 742 350 978 430
rect 1094 350 1482 430
rect 1598 350 1986 430
rect 2102 350 2490 430
rect 2606 350 2994 430
rect 3110 350 3498 430
rect 3614 350 4002 430
rect 4118 350 4506 430
rect 4622 350 5010 430
rect 5126 350 5514 430
rect 5630 350 6018 430
rect 6134 350 6522 430
rect 6638 350 7026 430
rect 7142 350 7530 430
rect 7646 350 8034 430
rect 8150 350 8538 430
rect 8654 350 9042 430
rect 9158 350 9546 430
rect 9662 350 10050 430
rect 10166 350 10554 430
rect 10670 350 11058 430
rect 11174 350 11562 430
rect 11678 350 12066 430
rect 12182 350 12570 430
rect 12686 350 13074 430
rect 13190 350 13578 430
rect 13694 350 14082 430
rect 14198 350 14586 430
rect 14702 350 15090 430
rect 15206 350 15594 430
rect 15710 350 16098 430
rect 16214 350 16602 430
rect 16718 350 17106 430
rect 17222 350 17610 430
rect 17726 350 18114 430
rect 18230 350 18618 430
rect 18734 350 19122 430
rect 19238 350 19626 430
rect 19742 350 20130 430
rect 20246 350 20634 430
rect 20750 350 21138 430
rect 21254 350 21642 430
rect 21758 350 22146 430
rect 22262 350 22650 430
rect 22766 350 23154 430
rect 23270 350 23658 430
rect 23774 350 24162 430
rect 24278 350 24666 430
rect 24782 350 25170 430
rect 25286 350 25674 430
rect 25790 350 26178 430
rect 26294 350 26682 430
rect 26798 350 27186 430
rect 27302 350 27690 430
rect 27806 350 28194 430
rect 28310 350 28698 430
rect 28814 350 29202 430
rect 29318 350 29706 430
rect 29822 350 30210 430
rect 30326 350 30714 430
rect 30830 350 31218 430
rect 31334 350 31722 430
rect 31838 350 32226 430
rect 32342 350 32730 430
rect 32846 350 33234 430
rect 33350 350 33738 430
rect 33854 350 34242 430
rect 34358 350 34746 430
rect 34862 350 35250 430
rect 35366 350 35754 430
rect 35870 350 36258 430
rect 36374 350 36762 430
rect 36878 350 37266 430
rect 37382 350 37770 430
rect 37886 350 38274 430
rect 38390 350 38778 430
rect 38894 350 39282 430
rect 39398 350 39786 430
rect 39902 350 40290 430
rect 40406 350 40794 430
rect 40910 350 41298 430
rect 41414 350 41802 430
rect 41918 350 42306 430
rect 42422 350 42810 430
rect 42926 350 43314 430
rect 43430 350 43818 430
rect 43934 350 44322 430
rect 44438 350 44826 430
rect 44942 350 45330 430
rect 45446 350 45834 430
rect 45950 350 46970 430
<< metal3 >>
rect 0 74088 400 74144
rect 0 73472 400 73528
rect 46600 73304 47000 73360
rect 0 72856 400 72912
rect 0 72240 400 72296
rect 46600 72184 47000 72240
rect 0 71624 400 71680
rect 0 71008 400 71064
rect 46600 71064 47000 71120
rect 0 70392 400 70448
rect 46600 69944 47000 70000
rect 0 69776 400 69832
rect 0 69160 400 69216
rect 46600 68824 47000 68880
rect 0 68544 400 68600
rect 0 67928 400 67984
rect 46600 67704 47000 67760
rect 0 67312 400 67368
rect 0 66696 400 66752
rect 46600 66584 47000 66640
rect 0 66080 400 66136
rect 0 65464 400 65520
rect 46600 65464 47000 65520
rect 0 64848 400 64904
rect 46600 64344 47000 64400
rect 0 64232 400 64288
rect 0 63616 400 63672
rect 46600 63224 47000 63280
rect 0 63000 400 63056
rect 0 62384 400 62440
rect 46600 62104 47000 62160
rect 0 61768 400 61824
rect 0 61152 400 61208
rect 46600 60984 47000 61040
rect 0 60536 400 60592
rect 0 59920 400 59976
rect 46600 59864 47000 59920
rect 0 59304 400 59360
rect 0 58688 400 58744
rect 46600 58744 47000 58800
rect 0 58072 400 58128
rect 46600 57624 47000 57680
rect 0 57456 400 57512
rect 0 56840 400 56896
rect 46600 56504 47000 56560
rect 0 56224 400 56280
rect 0 55608 400 55664
rect 46600 55384 47000 55440
rect 0 54992 400 55048
rect 0 54376 400 54432
rect 46600 54264 47000 54320
rect 0 53760 400 53816
rect 0 53144 400 53200
rect 46600 53144 47000 53200
rect 0 52528 400 52584
rect 46600 52024 47000 52080
rect 0 51912 400 51968
rect 0 51296 400 51352
rect 46600 50904 47000 50960
rect 0 50680 400 50736
rect 0 50064 400 50120
rect 46600 49784 47000 49840
rect 0 49448 400 49504
rect 0 48832 400 48888
rect 46600 48664 47000 48720
rect 0 48216 400 48272
rect 0 47600 400 47656
rect 46600 47544 47000 47600
rect 0 46984 400 47040
rect 0 46368 400 46424
rect 46600 46424 47000 46480
rect 0 45752 400 45808
rect 46600 45304 47000 45360
rect 0 45136 400 45192
rect 0 44520 400 44576
rect 46600 44184 47000 44240
rect 0 43904 400 43960
rect 0 43288 400 43344
rect 46600 43064 47000 43120
rect 0 42672 400 42728
rect 0 42056 400 42112
rect 46600 41944 47000 42000
rect 0 41440 400 41496
rect 0 40824 400 40880
rect 46600 40824 47000 40880
rect 0 40208 400 40264
rect 46600 39704 47000 39760
rect 0 39592 400 39648
rect 0 38976 400 39032
rect 46600 38584 47000 38640
rect 0 38360 400 38416
rect 0 37744 400 37800
rect 46600 37464 47000 37520
rect 0 37128 400 37184
rect 0 36512 400 36568
rect 46600 36344 47000 36400
rect 0 35896 400 35952
rect 0 35280 400 35336
rect 46600 35224 47000 35280
rect 0 34664 400 34720
rect 0 34048 400 34104
rect 46600 34104 47000 34160
rect 0 33432 400 33488
rect 46600 32984 47000 33040
rect 0 32816 400 32872
rect 0 32200 400 32256
rect 46600 31864 47000 31920
rect 0 31584 400 31640
rect 0 30968 400 31024
rect 46600 30744 47000 30800
rect 0 30352 400 30408
rect 0 29736 400 29792
rect 46600 29624 47000 29680
rect 0 29120 400 29176
rect 0 28504 400 28560
rect 46600 28504 47000 28560
rect 0 27888 400 27944
rect 46600 27384 47000 27440
rect 0 27272 400 27328
rect 0 26656 400 26712
rect 46600 26264 47000 26320
rect 0 26040 400 26096
rect 0 25424 400 25480
rect 46600 25144 47000 25200
rect 0 24808 400 24864
rect 0 24192 400 24248
rect 46600 24024 47000 24080
rect 0 23576 400 23632
rect 0 22960 400 23016
rect 46600 22904 47000 22960
rect 0 22344 400 22400
rect 0 21728 400 21784
rect 46600 21784 47000 21840
rect 0 21112 400 21168
rect 46600 20664 47000 20720
rect 0 20496 400 20552
rect 0 19880 400 19936
rect 46600 19544 47000 19600
rect 0 19264 400 19320
rect 0 18648 400 18704
rect 46600 18424 47000 18480
rect 0 18032 400 18088
rect 0 17416 400 17472
rect 46600 17304 47000 17360
rect 0 16800 400 16856
rect 0 16184 400 16240
rect 46600 16184 47000 16240
rect 0 15568 400 15624
rect 46600 15064 47000 15120
rect 0 14952 400 15008
rect 0 14336 400 14392
rect 46600 13944 47000 14000
rect 0 13720 400 13776
rect 0 13104 400 13160
rect 46600 12824 47000 12880
rect 0 12488 400 12544
rect 0 11872 400 11928
rect 46600 11704 47000 11760
rect 0 11256 400 11312
rect 0 10640 400 10696
rect 46600 10584 47000 10640
rect 0 10024 400 10080
rect 0 9408 400 9464
rect 46600 9464 47000 9520
rect 0 8792 400 8848
rect 46600 8344 47000 8400
rect 0 8176 400 8232
rect 0 7560 400 7616
rect 46600 7224 47000 7280
rect 0 6944 400 7000
rect 0 6328 400 6384
rect 46600 6104 47000 6160
rect 0 5712 400 5768
rect 0 5096 400 5152
rect 46600 4984 47000 5040
rect 0 4480 400 4536
rect 0 3864 400 3920
rect 46600 3864 47000 3920
rect 0 3248 400 3304
rect 46600 2744 47000 2800
rect 0 2632 400 2688
rect 0 2016 400 2072
rect 46600 1624 47000 1680
rect 0 1400 400 1456
rect 0 784 400 840
<< obsm3 >>
rect 350 74174 46919 74970
rect 430 74058 46919 74174
rect 350 73558 46919 74058
rect 430 73442 46919 73558
rect 350 73390 46919 73442
rect 350 73274 46570 73390
rect 350 72942 46919 73274
rect 430 72826 46919 72942
rect 350 72326 46919 72826
rect 430 72270 46919 72326
rect 430 72210 46570 72270
rect 350 72154 46570 72210
rect 350 71710 46919 72154
rect 430 71594 46919 71710
rect 350 71150 46919 71594
rect 350 71094 46570 71150
rect 430 71034 46570 71094
rect 430 70978 46919 71034
rect 350 70478 46919 70978
rect 430 70362 46919 70478
rect 350 70030 46919 70362
rect 350 69914 46570 70030
rect 350 69862 46919 69914
rect 430 69746 46919 69862
rect 350 69246 46919 69746
rect 430 69130 46919 69246
rect 350 68910 46919 69130
rect 350 68794 46570 68910
rect 350 68630 46919 68794
rect 430 68514 46919 68630
rect 350 68014 46919 68514
rect 430 67898 46919 68014
rect 350 67790 46919 67898
rect 350 67674 46570 67790
rect 350 67398 46919 67674
rect 430 67282 46919 67398
rect 350 66782 46919 67282
rect 430 66670 46919 66782
rect 430 66666 46570 66670
rect 350 66554 46570 66666
rect 350 66166 46919 66554
rect 430 66050 46919 66166
rect 350 65550 46919 66050
rect 430 65434 46570 65550
rect 350 64934 46919 65434
rect 430 64818 46919 64934
rect 350 64430 46919 64818
rect 350 64318 46570 64430
rect 430 64314 46570 64318
rect 430 64202 46919 64314
rect 350 63702 46919 64202
rect 430 63586 46919 63702
rect 350 63310 46919 63586
rect 350 63194 46570 63310
rect 350 63086 46919 63194
rect 430 62970 46919 63086
rect 350 62470 46919 62970
rect 430 62354 46919 62470
rect 350 62190 46919 62354
rect 350 62074 46570 62190
rect 350 61854 46919 62074
rect 430 61738 46919 61854
rect 350 61238 46919 61738
rect 430 61122 46919 61238
rect 350 61070 46919 61122
rect 350 60954 46570 61070
rect 350 60622 46919 60954
rect 430 60506 46919 60622
rect 350 60006 46919 60506
rect 430 59950 46919 60006
rect 430 59890 46570 59950
rect 350 59834 46570 59890
rect 350 59390 46919 59834
rect 430 59274 46919 59390
rect 350 58830 46919 59274
rect 350 58774 46570 58830
rect 430 58714 46570 58774
rect 430 58658 46919 58714
rect 350 58158 46919 58658
rect 430 58042 46919 58158
rect 350 57710 46919 58042
rect 350 57594 46570 57710
rect 350 57542 46919 57594
rect 430 57426 46919 57542
rect 350 56926 46919 57426
rect 430 56810 46919 56926
rect 350 56590 46919 56810
rect 350 56474 46570 56590
rect 350 56310 46919 56474
rect 430 56194 46919 56310
rect 350 55694 46919 56194
rect 430 55578 46919 55694
rect 350 55470 46919 55578
rect 350 55354 46570 55470
rect 350 55078 46919 55354
rect 430 54962 46919 55078
rect 350 54462 46919 54962
rect 430 54350 46919 54462
rect 430 54346 46570 54350
rect 350 54234 46570 54346
rect 350 53846 46919 54234
rect 430 53730 46919 53846
rect 350 53230 46919 53730
rect 430 53114 46570 53230
rect 350 52614 46919 53114
rect 430 52498 46919 52614
rect 350 52110 46919 52498
rect 350 51998 46570 52110
rect 430 51994 46570 51998
rect 430 51882 46919 51994
rect 350 51382 46919 51882
rect 430 51266 46919 51382
rect 350 50990 46919 51266
rect 350 50874 46570 50990
rect 350 50766 46919 50874
rect 430 50650 46919 50766
rect 350 50150 46919 50650
rect 430 50034 46919 50150
rect 350 49870 46919 50034
rect 350 49754 46570 49870
rect 350 49534 46919 49754
rect 430 49418 46919 49534
rect 350 48918 46919 49418
rect 430 48802 46919 48918
rect 350 48750 46919 48802
rect 350 48634 46570 48750
rect 350 48302 46919 48634
rect 430 48186 46919 48302
rect 350 47686 46919 48186
rect 430 47630 46919 47686
rect 430 47570 46570 47630
rect 350 47514 46570 47570
rect 350 47070 46919 47514
rect 430 46954 46919 47070
rect 350 46510 46919 46954
rect 350 46454 46570 46510
rect 430 46394 46570 46454
rect 430 46338 46919 46394
rect 350 45838 46919 46338
rect 430 45722 46919 45838
rect 350 45390 46919 45722
rect 350 45274 46570 45390
rect 350 45222 46919 45274
rect 430 45106 46919 45222
rect 350 44606 46919 45106
rect 430 44490 46919 44606
rect 350 44270 46919 44490
rect 350 44154 46570 44270
rect 350 43990 46919 44154
rect 430 43874 46919 43990
rect 350 43374 46919 43874
rect 430 43258 46919 43374
rect 350 43150 46919 43258
rect 350 43034 46570 43150
rect 350 42758 46919 43034
rect 430 42642 46919 42758
rect 350 42142 46919 42642
rect 430 42030 46919 42142
rect 430 42026 46570 42030
rect 350 41914 46570 42026
rect 350 41526 46919 41914
rect 430 41410 46919 41526
rect 350 40910 46919 41410
rect 430 40794 46570 40910
rect 350 40294 46919 40794
rect 430 40178 46919 40294
rect 350 39790 46919 40178
rect 350 39678 46570 39790
rect 430 39674 46570 39678
rect 430 39562 46919 39674
rect 350 39062 46919 39562
rect 430 38946 46919 39062
rect 350 38670 46919 38946
rect 350 38554 46570 38670
rect 350 38446 46919 38554
rect 430 38330 46919 38446
rect 350 37830 46919 38330
rect 430 37714 46919 37830
rect 350 37550 46919 37714
rect 350 37434 46570 37550
rect 350 37214 46919 37434
rect 430 37098 46919 37214
rect 350 36598 46919 37098
rect 430 36482 46919 36598
rect 350 36430 46919 36482
rect 350 36314 46570 36430
rect 350 35982 46919 36314
rect 430 35866 46919 35982
rect 350 35366 46919 35866
rect 430 35310 46919 35366
rect 430 35250 46570 35310
rect 350 35194 46570 35250
rect 350 34750 46919 35194
rect 430 34634 46919 34750
rect 350 34190 46919 34634
rect 350 34134 46570 34190
rect 430 34074 46570 34134
rect 430 34018 46919 34074
rect 350 33518 46919 34018
rect 430 33402 46919 33518
rect 350 33070 46919 33402
rect 350 32954 46570 33070
rect 350 32902 46919 32954
rect 430 32786 46919 32902
rect 350 32286 46919 32786
rect 430 32170 46919 32286
rect 350 31950 46919 32170
rect 350 31834 46570 31950
rect 350 31670 46919 31834
rect 430 31554 46919 31670
rect 350 31054 46919 31554
rect 430 30938 46919 31054
rect 350 30830 46919 30938
rect 350 30714 46570 30830
rect 350 30438 46919 30714
rect 430 30322 46919 30438
rect 350 29822 46919 30322
rect 430 29710 46919 29822
rect 430 29706 46570 29710
rect 350 29594 46570 29706
rect 350 29206 46919 29594
rect 430 29090 46919 29206
rect 350 28590 46919 29090
rect 430 28474 46570 28590
rect 350 27974 46919 28474
rect 430 27858 46919 27974
rect 350 27470 46919 27858
rect 350 27358 46570 27470
rect 430 27354 46570 27358
rect 430 27242 46919 27354
rect 350 26742 46919 27242
rect 430 26626 46919 26742
rect 350 26350 46919 26626
rect 350 26234 46570 26350
rect 350 26126 46919 26234
rect 430 26010 46919 26126
rect 350 25510 46919 26010
rect 430 25394 46919 25510
rect 350 25230 46919 25394
rect 350 25114 46570 25230
rect 350 24894 46919 25114
rect 430 24778 46919 24894
rect 350 24278 46919 24778
rect 430 24162 46919 24278
rect 350 24110 46919 24162
rect 350 23994 46570 24110
rect 350 23662 46919 23994
rect 430 23546 46919 23662
rect 350 23046 46919 23546
rect 430 22990 46919 23046
rect 430 22930 46570 22990
rect 350 22874 46570 22930
rect 350 22430 46919 22874
rect 430 22314 46919 22430
rect 350 21870 46919 22314
rect 350 21814 46570 21870
rect 430 21754 46570 21814
rect 430 21698 46919 21754
rect 350 21198 46919 21698
rect 430 21082 46919 21198
rect 350 20750 46919 21082
rect 350 20634 46570 20750
rect 350 20582 46919 20634
rect 430 20466 46919 20582
rect 350 19966 46919 20466
rect 430 19850 46919 19966
rect 350 19630 46919 19850
rect 350 19514 46570 19630
rect 350 19350 46919 19514
rect 430 19234 46919 19350
rect 350 18734 46919 19234
rect 430 18618 46919 18734
rect 350 18510 46919 18618
rect 350 18394 46570 18510
rect 350 18118 46919 18394
rect 430 18002 46919 18118
rect 350 17502 46919 18002
rect 430 17390 46919 17502
rect 430 17386 46570 17390
rect 350 17274 46570 17386
rect 350 16886 46919 17274
rect 430 16770 46919 16886
rect 350 16270 46919 16770
rect 430 16154 46570 16270
rect 350 15654 46919 16154
rect 430 15538 46919 15654
rect 350 15150 46919 15538
rect 350 15038 46570 15150
rect 430 15034 46570 15038
rect 430 14922 46919 15034
rect 350 14422 46919 14922
rect 430 14306 46919 14422
rect 350 14030 46919 14306
rect 350 13914 46570 14030
rect 350 13806 46919 13914
rect 430 13690 46919 13806
rect 350 13190 46919 13690
rect 430 13074 46919 13190
rect 350 12910 46919 13074
rect 350 12794 46570 12910
rect 350 12574 46919 12794
rect 430 12458 46919 12574
rect 350 11958 46919 12458
rect 430 11842 46919 11958
rect 350 11790 46919 11842
rect 350 11674 46570 11790
rect 350 11342 46919 11674
rect 430 11226 46919 11342
rect 350 10726 46919 11226
rect 430 10670 46919 10726
rect 430 10610 46570 10670
rect 350 10554 46570 10610
rect 350 10110 46919 10554
rect 430 9994 46919 10110
rect 350 9550 46919 9994
rect 350 9494 46570 9550
rect 430 9434 46570 9494
rect 430 9378 46919 9434
rect 350 8878 46919 9378
rect 430 8762 46919 8878
rect 350 8430 46919 8762
rect 350 8314 46570 8430
rect 350 8262 46919 8314
rect 430 8146 46919 8262
rect 350 7646 46919 8146
rect 430 7530 46919 7646
rect 350 7310 46919 7530
rect 350 7194 46570 7310
rect 350 7030 46919 7194
rect 430 6914 46919 7030
rect 350 6414 46919 6914
rect 430 6298 46919 6414
rect 350 6190 46919 6298
rect 350 6074 46570 6190
rect 350 5798 46919 6074
rect 430 5682 46919 5798
rect 350 5182 46919 5682
rect 430 5070 46919 5182
rect 430 5066 46570 5070
rect 350 4954 46570 5066
rect 350 4566 46919 4954
rect 430 4450 46919 4566
rect 350 3950 46919 4450
rect 430 3834 46570 3950
rect 350 3334 46919 3834
rect 430 3218 46919 3334
rect 350 2830 46919 3218
rect 350 2718 46570 2830
rect 430 2714 46570 2718
rect 430 2602 46919 2714
rect 350 2102 46919 2602
rect 430 1986 46919 2102
rect 350 1710 46919 1986
rect 350 1594 46570 1710
rect 350 1486 46919 1594
rect 430 1370 46919 1486
rect 350 870 46919 1370
rect 430 798 46919 870
<< metal4 >>
rect 2224 1538 2384 73334
rect 2554 1538 2714 73334
rect 9904 1538 10064 73334
rect 10234 1538 10394 73334
rect 17584 1538 17744 73334
rect 17914 1538 18074 73334
rect 25264 1538 25424 73334
rect 25594 1538 25754 73334
rect 32944 1538 33104 73334
rect 33274 1538 33434 73334
rect 40624 1538 40784 73334
rect 40954 1538 41114 73334
<< obsm4 >>
rect 518 73364 46298 74639
rect 518 1689 2194 73364
rect 2414 1689 2524 73364
rect 2744 1689 9874 73364
rect 10094 1689 10204 73364
rect 10424 1689 17554 73364
rect 17774 1689 17884 73364
rect 18104 1689 25234 73364
rect 25454 1689 25564 73364
rect 25784 1689 32914 73364
rect 33134 1689 33244 73364
rect 33464 1689 40594 73364
rect 40814 1689 40924 73364
rect 41144 1689 46298 73364
<< metal5 >>
rect 642 69599 46342 69759
rect 642 65689 46342 65849
rect 642 61779 46342 61939
rect 642 57869 46342 58029
rect 642 53959 46342 54119
rect 642 50049 46342 50209
rect 642 46139 46342 46299
rect 642 42229 46342 42389
rect 642 38319 46342 38479
rect 642 34409 46342 34569
rect 642 30499 46342 30659
rect 642 26589 46342 26749
rect 642 22679 46342 22839
rect 642 18769 46342 18929
rect 642 14859 46342 15019
rect 642 10949 46342 11109
rect 642 7039 46342 7199
rect 642 3129 46342 3289
<< obsm5 >>
rect 510 69809 46306 73970
rect 510 69549 592 69809
rect 510 65899 46306 69549
rect 510 65639 592 65899
rect 510 61989 46306 65639
rect 510 61729 592 61989
rect 510 58079 46306 61729
rect 510 57819 592 58079
rect 510 54169 46306 57819
rect 510 53909 592 54169
rect 510 50259 46306 53909
rect 510 49999 592 50259
rect 510 46349 46306 49999
rect 510 46089 592 46349
rect 510 42439 46306 46089
rect 510 42179 592 42439
rect 510 38529 46306 42179
rect 510 38269 592 38529
rect 510 34619 46306 38269
rect 510 34359 592 34619
rect 510 30709 46306 34359
rect 510 30449 592 30709
rect 510 26799 46306 30449
rect 510 26539 592 26799
rect 510 22889 46306 26539
rect 510 22629 592 22889
rect 510 18979 46306 22629
rect 510 18719 592 18979
rect 510 15069 46306 18719
rect 510 14809 592 15069
rect 510 11159 46306 14809
rect 510 10899 592 11159
rect 510 7249 46306 10899
rect 510 6989 592 7249
rect 510 3339 46306 6989
rect 510 3079 592 3339
rect 510 1686 46306 3079
<< labels >>
rlabel metal4 s 2224 1538 2384 73334 6 VDD
port 1 nsew power bidirectional
rlabel metal4 s 9904 1538 10064 73334 6 VDD
port 1 nsew power bidirectional
rlabel metal4 s 17584 1538 17744 73334 6 VDD
port 1 nsew power bidirectional
rlabel metal4 s 25264 1538 25424 73334 6 VDD
port 1 nsew power bidirectional
rlabel metal4 s 32944 1538 33104 73334 6 VDD
port 1 nsew power bidirectional
rlabel metal4 s 40624 1538 40784 73334 6 VDD
port 1 nsew power bidirectional
rlabel metal5 s 642 3129 46342 3289 6 VDD
port 1 nsew power bidirectional
rlabel metal5 s 642 10949 46342 11109 6 VDD
port 1 nsew power bidirectional
rlabel metal5 s 642 18769 46342 18929 6 VDD
port 1 nsew power bidirectional
rlabel metal5 s 642 26589 46342 26749 6 VDD
port 1 nsew power bidirectional
rlabel metal5 s 642 34409 46342 34569 6 VDD
port 1 nsew power bidirectional
rlabel metal5 s 642 42229 46342 42389 6 VDD
port 1 nsew power bidirectional
rlabel metal5 s 642 50049 46342 50209 6 VDD
port 1 nsew power bidirectional
rlabel metal5 s 642 57869 46342 58029 6 VDD
port 1 nsew power bidirectional
rlabel metal5 s 642 65689 46342 65849 6 VDD
port 1 nsew power bidirectional
rlabel metal4 s 2554 1538 2714 73334 6 VSS
port 2 nsew ground bidirectional
rlabel metal4 s 10234 1538 10394 73334 6 VSS
port 2 nsew ground bidirectional
rlabel metal4 s 17914 1538 18074 73334 6 VSS
port 2 nsew ground bidirectional
rlabel metal4 s 25594 1538 25754 73334 6 VSS
port 2 nsew ground bidirectional
rlabel metal4 s 33274 1538 33434 73334 6 VSS
port 2 nsew ground bidirectional
rlabel metal4 s 40954 1538 41114 73334 6 VSS
port 2 nsew ground bidirectional
rlabel metal5 s 642 7039 46342 7199 6 VSS
port 2 nsew ground bidirectional
rlabel metal5 s 642 14859 46342 15019 6 VSS
port 2 nsew ground bidirectional
rlabel metal5 s 642 22679 46342 22839 6 VSS
port 2 nsew ground bidirectional
rlabel metal5 s 642 30499 46342 30659 6 VSS
port 2 nsew ground bidirectional
rlabel metal5 s 642 38319 46342 38479 6 VSS
port 2 nsew ground bidirectional
rlabel metal5 s 642 46139 46342 46299 6 VSS
port 2 nsew ground bidirectional
rlabel metal5 s 642 53959 46342 54119 6 VSS
port 2 nsew ground bidirectional
rlabel metal5 s 642 61779 46342 61939 6 VSS
port 2 nsew ground bidirectional
rlabel metal5 s 642 69599 46342 69759 6 VSS
port 2 nsew ground bidirectional
rlabel metal3 s 0 784 400 840 6 debug_in
port 3 nsew signal output
rlabel metal3 s 0 1400 400 1456 6 debug_mode
port 4 nsew signal input
rlabel metal3 s 0 2016 400 2072 6 debug_oeb
port 5 nsew signal input
rlabel metal3 s 0 2632 400 2688 6 debug_out
port 6 nsew signal input
rlabel metal3 s 0 3864 400 3920 6 irq[0]
port 7 nsew signal output
rlabel metal3 s 0 4480 400 4536 6 irq[1]
port 8 nsew signal output
rlabel metal3 s 0 5096 400 5152 6 irq[2]
port 9 nsew signal output
rlabel metal2 s 29736 0 29792 400 6 mask_rev_in[0]
port 10 nsew signal input
rlabel metal2 s 34776 0 34832 400 6 mask_rev_in[10]
port 11 nsew signal input
rlabel metal2 s 35280 0 35336 400 6 mask_rev_in[11]
port 12 nsew signal input
rlabel metal2 s 35784 0 35840 400 6 mask_rev_in[12]
port 13 nsew signal input
rlabel metal2 s 36288 0 36344 400 6 mask_rev_in[13]
port 14 nsew signal input
rlabel metal2 s 36792 0 36848 400 6 mask_rev_in[14]
port 15 nsew signal input
rlabel metal2 s 37296 0 37352 400 6 mask_rev_in[15]
port 16 nsew signal input
rlabel metal2 s 37800 0 37856 400 6 mask_rev_in[16]
port 17 nsew signal input
rlabel metal2 s 38304 0 38360 400 6 mask_rev_in[17]
port 18 nsew signal input
rlabel metal2 s 38808 0 38864 400 6 mask_rev_in[18]
port 19 nsew signal input
rlabel metal2 s 39312 0 39368 400 6 mask_rev_in[19]
port 20 nsew signal input
rlabel metal2 s 30240 0 30296 400 6 mask_rev_in[1]
port 21 nsew signal input
rlabel metal2 s 39816 0 39872 400 6 mask_rev_in[20]
port 22 nsew signal input
rlabel metal2 s 40320 0 40376 400 6 mask_rev_in[21]
port 23 nsew signal input
rlabel metal2 s 40824 0 40880 400 6 mask_rev_in[22]
port 24 nsew signal input
rlabel metal2 s 41328 0 41384 400 6 mask_rev_in[23]
port 25 nsew signal input
rlabel metal2 s 41832 0 41888 400 6 mask_rev_in[24]
port 26 nsew signal input
rlabel metal2 s 42336 0 42392 400 6 mask_rev_in[25]
port 27 nsew signal input
rlabel metal2 s 42840 0 42896 400 6 mask_rev_in[26]
port 28 nsew signal input
rlabel metal2 s 43344 0 43400 400 6 mask_rev_in[27]
port 29 nsew signal input
rlabel metal2 s 43848 0 43904 400 6 mask_rev_in[28]
port 30 nsew signal input
rlabel metal2 s 44352 0 44408 400 6 mask_rev_in[29]
port 31 nsew signal input
rlabel metal2 s 30744 0 30800 400 6 mask_rev_in[2]
port 32 nsew signal input
rlabel metal2 s 44856 0 44912 400 6 mask_rev_in[30]
port 33 nsew signal input
rlabel metal2 s 45360 0 45416 400 6 mask_rev_in[31]
port 34 nsew signal input
rlabel metal2 s 31248 0 31304 400 6 mask_rev_in[3]
port 35 nsew signal input
rlabel metal2 s 31752 0 31808 400 6 mask_rev_in[4]
port 36 nsew signal input
rlabel metal2 s 32256 0 32312 400 6 mask_rev_in[5]
port 37 nsew signal input
rlabel metal2 s 32760 0 32816 400 6 mask_rev_in[6]
port 38 nsew signal input
rlabel metal2 s 33264 0 33320 400 6 mask_rev_in[7]
port 39 nsew signal input
rlabel metal2 s 33768 0 33824 400 6 mask_rev_in[8]
port 40 nsew signal input
rlabel metal2 s 34272 0 34328 400 6 mask_rev_in[9]
port 41 nsew signal input
rlabel metal3 s 46600 7224 47000 7280 6 mgmt_gpio_in[0]
port 42 nsew signal input
rlabel metal3 s 46600 40824 47000 40880 6 mgmt_gpio_in[10]
port 43 nsew signal input
rlabel metal3 s 46600 44184 47000 44240 6 mgmt_gpio_in[11]
port 44 nsew signal input
rlabel metal3 s 46600 47544 47000 47600 6 mgmt_gpio_in[12]
port 45 nsew signal input
rlabel metal3 s 46600 50904 47000 50960 6 mgmt_gpio_in[13]
port 46 nsew signal input
rlabel metal3 s 46600 54264 47000 54320 6 mgmt_gpio_in[14]
port 47 nsew signal input
rlabel metal3 s 46600 57624 47000 57680 6 mgmt_gpio_in[15]
port 48 nsew signal input
rlabel metal3 s 46600 60984 47000 61040 6 mgmt_gpio_in[16]
port 49 nsew signal input
rlabel metal3 s 46600 64344 47000 64400 6 mgmt_gpio_in[17]
port 50 nsew signal input
rlabel metal3 s 46600 67704 47000 67760 6 mgmt_gpio_in[18]
port 51 nsew signal input
rlabel metal3 s 46600 71064 47000 71120 6 mgmt_gpio_in[19]
port 52 nsew signal input
rlabel metal3 s 46600 10584 47000 10640 6 mgmt_gpio_in[1]
port 53 nsew signal input
rlabel metal3 s 0 41440 400 41496 6 mgmt_gpio_in[20]
port 54 nsew signal input
rlabel metal3 s 0 43288 400 43344 6 mgmt_gpio_in[21]
port 55 nsew signal input
rlabel metal3 s 0 45136 400 45192 6 mgmt_gpio_in[22]
port 56 nsew signal input
rlabel metal3 s 0 46984 400 47040 6 mgmt_gpio_in[23]
port 57 nsew signal input
rlabel metal3 s 0 48832 400 48888 6 mgmt_gpio_in[24]
port 58 nsew signal input
rlabel metal3 s 0 50680 400 50736 6 mgmt_gpio_in[25]
port 59 nsew signal input
rlabel metal3 s 0 52528 400 52584 6 mgmt_gpio_in[26]
port 60 nsew signal input
rlabel metal3 s 0 54376 400 54432 6 mgmt_gpio_in[27]
port 61 nsew signal input
rlabel metal3 s 0 56224 400 56280 6 mgmt_gpio_in[28]
port 62 nsew signal input
rlabel metal3 s 0 58072 400 58128 6 mgmt_gpio_in[29]
port 63 nsew signal input
rlabel metal3 s 46600 13944 47000 14000 6 mgmt_gpio_in[2]
port 64 nsew signal input
rlabel metal3 s 0 59920 400 59976 6 mgmt_gpio_in[30]
port 65 nsew signal input
rlabel metal3 s 0 61768 400 61824 6 mgmt_gpio_in[31]
port 66 nsew signal input
rlabel metal3 s 0 63616 400 63672 6 mgmt_gpio_in[32]
port 67 nsew signal input
rlabel metal3 s 0 65464 400 65520 6 mgmt_gpio_in[33]
port 68 nsew signal input
rlabel metal3 s 0 67312 400 67368 6 mgmt_gpio_in[34]
port 69 nsew signal input
rlabel metal3 s 0 69160 400 69216 6 mgmt_gpio_in[35]
port 70 nsew signal input
rlabel metal3 s 0 71008 400 71064 6 mgmt_gpio_in[36]
port 71 nsew signal input
rlabel metal3 s 0 72856 400 72912 6 mgmt_gpio_in[37]
port 72 nsew signal input
rlabel metal3 s 46600 17304 47000 17360 6 mgmt_gpio_in[3]
port 73 nsew signal input
rlabel metal3 s 46600 20664 47000 20720 6 mgmt_gpio_in[4]
port 74 nsew signal input
rlabel metal3 s 46600 24024 47000 24080 6 mgmt_gpio_in[5]
port 75 nsew signal input
rlabel metal3 s 46600 27384 47000 27440 6 mgmt_gpio_in[6]
port 76 nsew signal input
rlabel metal3 s 46600 30744 47000 30800 6 mgmt_gpio_in[7]
port 77 nsew signal input
rlabel metal3 s 46600 34104 47000 34160 6 mgmt_gpio_in[8]
port 78 nsew signal input
rlabel metal3 s 46600 37464 47000 37520 6 mgmt_gpio_in[9]
port 79 nsew signal input
rlabel metal3 s 46600 8344 47000 8400 6 mgmt_gpio_oeb[0]
port 80 nsew signal output
rlabel metal3 s 46600 41944 47000 42000 6 mgmt_gpio_oeb[10]
port 81 nsew signal output
rlabel metal3 s 46600 45304 47000 45360 6 mgmt_gpio_oeb[11]
port 82 nsew signal output
rlabel metal3 s 46600 48664 47000 48720 6 mgmt_gpio_oeb[12]
port 83 nsew signal output
rlabel metal3 s 46600 52024 47000 52080 6 mgmt_gpio_oeb[13]
port 84 nsew signal output
rlabel metal3 s 46600 55384 47000 55440 6 mgmt_gpio_oeb[14]
port 85 nsew signal output
rlabel metal3 s 46600 58744 47000 58800 6 mgmt_gpio_oeb[15]
port 86 nsew signal output
rlabel metal3 s 46600 62104 47000 62160 6 mgmt_gpio_oeb[16]
port 87 nsew signal output
rlabel metal3 s 46600 65464 47000 65520 6 mgmt_gpio_oeb[17]
port 88 nsew signal output
rlabel metal3 s 46600 68824 47000 68880 6 mgmt_gpio_oeb[18]
port 89 nsew signal output
rlabel metal3 s 46600 72184 47000 72240 6 mgmt_gpio_oeb[19]
port 90 nsew signal output
rlabel metal3 s 46600 11704 47000 11760 6 mgmt_gpio_oeb[1]
port 91 nsew signal output
rlabel metal3 s 0 42056 400 42112 6 mgmt_gpio_oeb[20]
port 92 nsew signal output
rlabel metal3 s 0 43904 400 43960 6 mgmt_gpio_oeb[21]
port 93 nsew signal output
rlabel metal3 s 0 45752 400 45808 6 mgmt_gpio_oeb[22]
port 94 nsew signal output
rlabel metal3 s 0 47600 400 47656 6 mgmt_gpio_oeb[23]
port 95 nsew signal output
rlabel metal3 s 0 49448 400 49504 6 mgmt_gpio_oeb[24]
port 96 nsew signal output
rlabel metal3 s 0 51296 400 51352 6 mgmt_gpio_oeb[25]
port 97 nsew signal output
rlabel metal3 s 0 53144 400 53200 6 mgmt_gpio_oeb[26]
port 98 nsew signal output
rlabel metal3 s 0 54992 400 55048 6 mgmt_gpio_oeb[27]
port 99 nsew signal output
rlabel metal3 s 0 56840 400 56896 6 mgmt_gpio_oeb[28]
port 100 nsew signal output
rlabel metal3 s 0 58688 400 58744 6 mgmt_gpio_oeb[29]
port 101 nsew signal output
rlabel metal3 s 46600 15064 47000 15120 6 mgmt_gpio_oeb[2]
port 102 nsew signal output
rlabel metal3 s 0 60536 400 60592 6 mgmt_gpio_oeb[30]
port 103 nsew signal output
rlabel metal3 s 0 62384 400 62440 6 mgmt_gpio_oeb[31]
port 104 nsew signal output
rlabel metal3 s 0 64232 400 64288 6 mgmt_gpio_oeb[32]
port 105 nsew signal output
rlabel metal3 s 0 66080 400 66136 6 mgmt_gpio_oeb[33]
port 106 nsew signal output
rlabel metal3 s 0 67928 400 67984 6 mgmt_gpio_oeb[34]
port 107 nsew signal output
rlabel metal3 s 0 69776 400 69832 6 mgmt_gpio_oeb[35]
port 108 nsew signal output
rlabel metal3 s 0 71624 400 71680 6 mgmt_gpio_oeb[36]
port 109 nsew signal output
rlabel metal3 s 0 73472 400 73528 6 mgmt_gpio_oeb[37]
port 110 nsew signal output
rlabel metal3 s 46600 18424 47000 18480 6 mgmt_gpio_oeb[3]
port 111 nsew signal output
rlabel metal3 s 46600 21784 47000 21840 6 mgmt_gpio_oeb[4]
port 112 nsew signal output
rlabel metal3 s 46600 25144 47000 25200 6 mgmt_gpio_oeb[5]
port 113 nsew signal output
rlabel metal3 s 46600 28504 47000 28560 6 mgmt_gpio_oeb[6]
port 114 nsew signal output
rlabel metal3 s 46600 31864 47000 31920 6 mgmt_gpio_oeb[7]
port 115 nsew signal output
rlabel metal3 s 46600 35224 47000 35280 6 mgmt_gpio_oeb[8]
port 116 nsew signal output
rlabel metal3 s 46600 38584 47000 38640 6 mgmt_gpio_oeb[9]
port 117 nsew signal output
rlabel metal3 s 46600 9464 47000 9520 6 mgmt_gpio_out[0]
port 118 nsew signal output
rlabel metal3 s 46600 43064 47000 43120 6 mgmt_gpio_out[10]
port 119 nsew signal output
rlabel metal3 s 46600 46424 47000 46480 6 mgmt_gpio_out[11]
port 120 nsew signal output
rlabel metal3 s 46600 49784 47000 49840 6 mgmt_gpio_out[12]
port 121 nsew signal output
rlabel metal3 s 46600 53144 47000 53200 6 mgmt_gpio_out[13]
port 122 nsew signal output
rlabel metal3 s 46600 56504 47000 56560 6 mgmt_gpio_out[14]
port 123 nsew signal output
rlabel metal3 s 46600 59864 47000 59920 6 mgmt_gpio_out[15]
port 124 nsew signal output
rlabel metal3 s 46600 63224 47000 63280 6 mgmt_gpio_out[16]
port 125 nsew signal output
rlabel metal3 s 46600 66584 47000 66640 6 mgmt_gpio_out[17]
port 126 nsew signal output
rlabel metal3 s 46600 69944 47000 70000 6 mgmt_gpio_out[18]
port 127 nsew signal output
rlabel metal3 s 46600 73304 47000 73360 6 mgmt_gpio_out[19]
port 128 nsew signal output
rlabel metal3 s 46600 12824 47000 12880 6 mgmt_gpio_out[1]
port 129 nsew signal output
rlabel metal3 s 0 42672 400 42728 6 mgmt_gpio_out[20]
port 130 nsew signal output
rlabel metal3 s 0 44520 400 44576 6 mgmt_gpio_out[21]
port 131 nsew signal output
rlabel metal3 s 0 46368 400 46424 6 mgmt_gpio_out[22]
port 132 nsew signal output
rlabel metal3 s 0 48216 400 48272 6 mgmt_gpio_out[23]
port 133 nsew signal output
rlabel metal3 s 0 50064 400 50120 6 mgmt_gpio_out[24]
port 134 nsew signal output
rlabel metal3 s 0 51912 400 51968 6 mgmt_gpio_out[25]
port 135 nsew signal output
rlabel metal3 s 0 53760 400 53816 6 mgmt_gpio_out[26]
port 136 nsew signal output
rlabel metal3 s 0 55608 400 55664 6 mgmt_gpio_out[27]
port 137 nsew signal output
rlabel metal3 s 0 57456 400 57512 6 mgmt_gpio_out[28]
port 138 nsew signal output
rlabel metal3 s 0 59304 400 59360 6 mgmt_gpio_out[29]
port 139 nsew signal output
rlabel metal3 s 46600 16184 47000 16240 6 mgmt_gpio_out[2]
port 140 nsew signal output
rlabel metal3 s 0 61152 400 61208 6 mgmt_gpio_out[30]
port 141 nsew signal output
rlabel metal3 s 0 63000 400 63056 6 mgmt_gpio_out[31]
port 142 nsew signal output
rlabel metal3 s 0 64848 400 64904 6 mgmt_gpio_out[32]
port 143 nsew signal output
rlabel metal3 s 0 66696 400 66752 6 mgmt_gpio_out[33]
port 144 nsew signal output
rlabel metal3 s 0 68544 400 68600 6 mgmt_gpio_out[34]
port 145 nsew signal output
rlabel metal3 s 0 70392 400 70448 6 mgmt_gpio_out[35]
port 146 nsew signal output
rlabel metal3 s 0 72240 400 72296 6 mgmt_gpio_out[36]
port 147 nsew signal output
rlabel metal3 s 0 74088 400 74144 6 mgmt_gpio_out[37]
port 148 nsew signal output
rlabel metal3 s 46600 19544 47000 19600 6 mgmt_gpio_out[3]
port 149 nsew signal output
rlabel metal3 s 46600 22904 47000 22960 6 mgmt_gpio_out[4]
port 150 nsew signal output
rlabel metal3 s 46600 26264 47000 26320 6 mgmt_gpio_out[5]
port 151 nsew signal output
rlabel metal3 s 46600 29624 47000 29680 6 mgmt_gpio_out[6]
port 152 nsew signal output
rlabel metal3 s 46600 32984 47000 33040 6 mgmt_gpio_out[7]
port 153 nsew signal output
rlabel metal3 s 46600 36344 47000 36400 6 mgmt_gpio_out[8]
port 154 nsew signal output
rlabel metal3 s 46600 39704 47000 39760 6 mgmt_gpio_out[9]
port 155 nsew signal output
rlabel metal2 s 1512 0 1568 400 6 pad_flash_clk
port 156 nsew signal output
rlabel metal2 s 2016 0 2072 400 6 pad_flash_clk_oe
port 157 nsew signal output
rlabel metal2 s 2520 0 2576 400 6 pad_flash_csb
port 158 nsew signal output
rlabel metal2 s 3024 0 3080 400 6 pad_flash_csb_oe
port 159 nsew signal output
rlabel metal2 s 3528 0 3584 400 6 pad_flash_io0_di
port 160 nsew signal input
rlabel metal2 s 4032 0 4088 400 6 pad_flash_io0_do
port 161 nsew signal output
rlabel metal2 s 4536 0 4592 400 6 pad_flash_io0_ie
port 162 nsew signal output
rlabel metal2 s 5040 0 5096 400 6 pad_flash_io0_oe
port 163 nsew signal output
rlabel metal2 s 5544 0 5600 400 6 pad_flash_io1_di
port 164 nsew signal input
rlabel metal2 s 6048 0 6104 400 6 pad_flash_io1_do
port 165 nsew signal output
rlabel metal2 s 6552 0 6608 400 6 pad_flash_io1_ie
port 166 nsew signal output
rlabel metal2 s 7056 0 7112 400 6 pad_flash_io1_oe
port 167 nsew signal output
rlabel metal2 s 13608 0 13664 400 6 pll90_sel[0]
port 168 nsew signal output
rlabel metal2 s 14112 0 14168 400 6 pll90_sel[1]
port 169 nsew signal output
rlabel metal2 s 14616 0 14672 400 6 pll90_sel[2]
port 170 nsew signal output
rlabel metal2 s 28224 0 28280 400 6 pll_bypass
port 171 nsew signal output
rlabel metal2 s 9072 0 9128 400 6 pll_dco_ena
port 172 nsew signal output
rlabel metal2 s 9576 0 9632 400 6 pll_div[0]
port 173 nsew signal output
rlabel metal2 s 10080 0 10136 400 6 pll_div[1]
port 174 nsew signal output
rlabel metal2 s 10584 0 10640 400 6 pll_div[2]
port 175 nsew signal output
rlabel metal2 s 11088 0 11144 400 6 pll_div[3]
port 176 nsew signal output
rlabel metal2 s 11592 0 11648 400 6 pll_div[4]
port 177 nsew signal output
rlabel metal2 s 8568 0 8624 400 6 pll_ena
port 178 nsew signal output
rlabel metal2 s 12096 0 12152 400 6 pll_sel[0]
port 179 nsew signal output
rlabel metal2 s 12600 0 12656 400 6 pll_sel[1]
port 180 nsew signal output
rlabel metal2 s 13104 0 13160 400 6 pll_sel[2]
port 181 nsew signal output
rlabel metal2 s 15120 0 15176 400 6 pll_trim[0]
port 182 nsew signal output
rlabel metal2 s 20160 0 20216 400 6 pll_trim[10]
port 183 nsew signal output
rlabel metal2 s 20664 0 20720 400 6 pll_trim[11]
port 184 nsew signal output
rlabel metal2 s 21168 0 21224 400 6 pll_trim[12]
port 185 nsew signal output
rlabel metal2 s 21672 0 21728 400 6 pll_trim[13]
port 186 nsew signal output
rlabel metal2 s 22176 0 22232 400 6 pll_trim[14]
port 187 nsew signal output
rlabel metal2 s 22680 0 22736 400 6 pll_trim[15]
port 188 nsew signal output
rlabel metal2 s 23184 0 23240 400 6 pll_trim[16]
port 189 nsew signal output
rlabel metal2 s 23688 0 23744 400 6 pll_trim[17]
port 190 nsew signal output
rlabel metal2 s 24192 0 24248 400 6 pll_trim[18]
port 191 nsew signal output
rlabel metal2 s 24696 0 24752 400 6 pll_trim[19]
port 192 nsew signal output
rlabel metal2 s 15624 0 15680 400 6 pll_trim[1]
port 193 nsew signal output
rlabel metal2 s 25200 0 25256 400 6 pll_trim[20]
port 194 nsew signal output
rlabel metal2 s 25704 0 25760 400 6 pll_trim[21]
port 195 nsew signal output
rlabel metal2 s 26208 0 26264 400 6 pll_trim[22]
port 196 nsew signal output
rlabel metal2 s 26712 0 26768 400 6 pll_trim[23]
port 197 nsew signal output
rlabel metal2 s 27216 0 27272 400 6 pll_trim[24]
port 198 nsew signal output
rlabel metal2 s 27720 0 27776 400 6 pll_trim[25]
port 199 nsew signal output
rlabel metal2 s 16128 0 16184 400 6 pll_trim[2]
port 200 nsew signal output
rlabel metal2 s 16632 0 16688 400 6 pll_trim[3]
port 201 nsew signal output
rlabel metal2 s 17136 0 17192 400 6 pll_trim[4]
port 202 nsew signal output
rlabel metal2 s 17640 0 17696 400 6 pll_trim[5]
port 203 nsew signal output
rlabel metal2 s 18144 0 18200 400 6 pll_trim[6]
port 204 nsew signal output
rlabel metal2 s 18648 0 18704 400 6 pll_trim[7]
port 205 nsew signal output
rlabel metal2 s 19152 0 19208 400 6 pll_trim[8]
port 206 nsew signal output
rlabel metal2 s 19656 0 19712 400 6 pll_trim[9]
port 207 nsew signal output
rlabel metal2 s 7560 0 7616 400 6 porb
port 208 nsew signal input
rlabel metal2 s 45864 0 45920 400 6 pwr_ctrl_out
port 209 nsew signal output
rlabel metal3 s 0 10024 400 10080 6 qspi_enabled
port 210 nsew signal input
rlabel metal2 s 8064 0 8120 400 6 reset
port 211 nsew signal output
rlabel metal3 s 0 9408 400 9464 6 ser_rx
port 212 nsew signal output
rlabel metal3 s 0 8792 400 8848 6 ser_tx
port 213 nsew signal input
rlabel metal3 s 46600 1624 47000 1680 6 serial_clock
port 214 nsew signal output
rlabel metal3 s 46600 4984 47000 5040 6 serial_data_1
port 215 nsew signal output
rlabel metal3 s 46600 6104 47000 6160 6 serial_data_2
port 216 nsew signal output
rlabel metal3 s 46600 3864 47000 3920 6 serial_load
port 217 nsew signal output
rlabel metal3 s 46600 2744 47000 2800 6 serial_resetn
port 218 nsew signal output
rlabel metal3 s 0 7560 400 7616 6 spi_csb
port 219 nsew signal input
rlabel metal3 s 0 11256 400 11312 6 spi_enabled
port 220 nsew signal input
rlabel metal3 s 0 6944 400 7000 6 spi_sck
port 221 nsew signal input
rlabel metal3 s 0 8176 400 8232 6 spi_sdi
port 222 nsew signal output
rlabel metal3 s 0 6328 400 6384 6 spi_sdo
port 223 nsew signal input
rlabel metal3 s 0 5712 400 5768 6 spi_sdoenb
port 224 nsew signal input
rlabel metal3 s 0 32816 400 32872 6 spimemio_flash_clk
port 225 nsew signal input
rlabel metal3 s 0 33432 400 33488 6 spimemio_flash_csb
port 226 nsew signal input
rlabel metal3 s 0 34048 400 34104 6 spimemio_flash_io0_di
port 227 nsew signal output
rlabel metal3 s 0 34664 400 34720 6 spimemio_flash_io0_do
port 228 nsew signal input
rlabel metal3 s 0 35280 400 35336 6 spimemio_flash_io0_oeb
port 229 nsew signal input
rlabel metal3 s 0 35896 400 35952 6 spimemio_flash_io1_di
port 230 nsew signal output
rlabel metal3 s 0 36512 400 36568 6 spimemio_flash_io1_do
port 231 nsew signal input
rlabel metal3 s 0 37128 400 37184 6 spimemio_flash_io1_oeb
port 232 nsew signal input
rlabel metal3 s 0 37744 400 37800 6 spimemio_flash_io2_di
port 233 nsew signal output
rlabel metal3 s 0 38360 400 38416 6 spimemio_flash_io2_do
port 234 nsew signal input
rlabel metal3 s 0 38976 400 39032 6 spimemio_flash_io2_oeb
port 235 nsew signal input
rlabel metal3 s 0 39592 400 39648 6 spimemio_flash_io3_di
port 236 nsew signal output
rlabel metal3 s 0 40208 400 40264 6 spimemio_flash_io3_do
port 237 nsew signal input
rlabel metal3 s 0 40824 400 40880 6 spimemio_flash_io3_oeb
port 238 nsew signal input
rlabel metal3 s 0 3248 400 3304 6 trap
port 239 nsew signal input
rlabel metal3 s 0 10640 400 10696 6 uart_enabled
port 240 nsew signal input
rlabel metal2 s 1008 0 1064 400 6 user_clock
port 241 nsew signal input
rlabel metal3 s 0 11872 400 11928 6 wb_ack_o
port 242 nsew signal output
rlabel metal2 s 2184 74600 2240 75000 6 wb_adr_i[0]
port 243 nsew signal input
rlabel metal2 s 8344 74600 8400 75000 6 wb_adr_i[10]
port 244 nsew signal input
rlabel metal2 s 8960 74600 9016 75000 6 wb_adr_i[11]
port 245 nsew signal input
rlabel metal2 s 9576 74600 9632 75000 6 wb_adr_i[12]
port 246 nsew signal input
rlabel metal2 s 10192 74600 10248 75000 6 wb_adr_i[13]
port 247 nsew signal input
rlabel metal2 s 10808 74600 10864 75000 6 wb_adr_i[14]
port 248 nsew signal input
rlabel metal2 s 11424 74600 11480 75000 6 wb_adr_i[15]
port 249 nsew signal input
rlabel metal2 s 12040 74600 12096 75000 6 wb_adr_i[16]
port 250 nsew signal input
rlabel metal2 s 12656 74600 12712 75000 6 wb_adr_i[17]
port 251 nsew signal input
rlabel metal2 s 13272 74600 13328 75000 6 wb_adr_i[18]
port 252 nsew signal input
rlabel metal2 s 13888 74600 13944 75000 6 wb_adr_i[19]
port 253 nsew signal input
rlabel metal2 s 2800 74600 2856 75000 6 wb_adr_i[1]
port 254 nsew signal input
rlabel metal2 s 14504 74600 14560 75000 6 wb_adr_i[20]
port 255 nsew signal input
rlabel metal2 s 15120 74600 15176 75000 6 wb_adr_i[21]
port 256 nsew signal input
rlabel metal2 s 15736 74600 15792 75000 6 wb_adr_i[22]
port 257 nsew signal input
rlabel metal2 s 16352 74600 16408 75000 6 wb_adr_i[23]
port 258 nsew signal input
rlabel metal2 s 16968 74600 17024 75000 6 wb_adr_i[24]
port 259 nsew signal input
rlabel metal2 s 17584 74600 17640 75000 6 wb_adr_i[25]
port 260 nsew signal input
rlabel metal2 s 18200 74600 18256 75000 6 wb_adr_i[26]
port 261 nsew signal input
rlabel metal2 s 18816 74600 18872 75000 6 wb_adr_i[27]
port 262 nsew signal input
rlabel metal2 s 19432 74600 19488 75000 6 wb_adr_i[28]
port 263 nsew signal input
rlabel metal2 s 20048 74600 20104 75000 6 wb_adr_i[29]
port 264 nsew signal input
rlabel metal2 s 3416 74600 3472 75000 6 wb_adr_i[2]
port 265 nsew signal input
rlabel metal2 s 20664 74600 20720 75000 6 wb_adr_i[30]
port 266 nsew signal input
rlabel metal2 s 21280 74600 21336 75000 6 wb_adr_i[31]
port 267 nsew signal input
rlabel metal2 s 4032 74600 4088 75000 6 wb_adr_i[3]
port 268 nsew signal input
rlabel metal2 s 4648 74600 4704 75000 6 wb_adr_i[4]
port 269 nsew signal input
rlabel metal2 s 5264 74600 5320 75000 6 wb_adr_i[5]
port 270 nsew signal input
rlabel metal2 s 5880 74600 5936 75000 6 wb_adr_i[6]
port 271 nsew signal input
rlabel metal2 s 6496 74600 6552 75000 6 wb_adr_i[7]
port 272 nsew signal input
rlabel metal2 s 7112 74600 7168 75000 6 wb_adr_i[8]
port 273 nsew signal input
rlabel metal2 s 7728 74600 7784 75000 6 wb_adr_i[9]
port 274 nsew signal input
rlabel metal2 s 28728 0 28784 400 6 wb_clk_i
port 275 nsew signal input
rlabel metal2 s 44688 74600 44744 75000 6 wb_cyc_i
port 276 nsew signal input
rlabel metal2 s 21896 74600 21952 75000 6 wb_dat_i[0]
port 277 nsew signal input
rlabel metal2 s 28056 74600 28112 75000 6 wb_dat_i[10]
port 278 nsew signal input
rlabel metal2 s 28672 74600 28728 75000 6 wb_dat_i[11]
port 279 nsew signal input
rlabel metal2 s 29288 74600 29344 75000 6 wb_dat_i[12]
port 280 nsew signal input
rlabel metal2 s 29904 74600 29960 75000 6 wb_dat_i[13]
port 281 nsew signal input
rlabel metal2 s 30520 74600 30576 75000 6 wb_dat_i[14]
port 282 nsew signal input
rlabel metal2 s 31136 74600 31192 75000 6 wb_dat_i[15]
port 283 nsew signal input
rlabel metal2 s 31752 74600 31808 75000 6 wb_dat_i[16]
port 284 nsew signal input
rlabel metal2 s 32368 74600 32424 75000 6 wb_dat_i[17]
port 285 nsew signal input
rlabel metal2 s 32984 74600 33040 75000 6 wb_dat_i[18]
port 286 nsew signal input
rlabel metal2 s 33600 74600 33656 75000 6 wb_dat_i[19]
port 287 nsew signal input
rlabel metal2 s 22512 74600 22568 75000 6 wb_dat_i[1]
port 288 nsew signal input
rlabel metal2 s 34216 74600 34272 75000 6 wb_dat_i[20]
port 289 nsew signal input
rlabel metal2 s 34832 74600 34888 75000 6 wb_dat_i[21]
port 290 nsew signal input
rlabel metal2 s 35448 74600 35504 75000 6 wb_dat_i[22]
port 291 nsew signal input
rlabel metal2 s 36064 74600 36120 75000 6 wb_dat_i[23]
port 292 nsew signal input
rlabel metal2 s 36680 74600 36736 75000 6 wb_dat_i[24]
port 293 nsew signal input
rlabel metal2 s 37296 74600 37352 75000 6 wb_dat_i[25]
port 294 nsew signal input
rlabel metal2 s 37912 74600 37968 75000 6 wb_dat_i[26]
port 295 nsew signal input
rlabel metal2 s 38528 74600 38584 75000 6 wb_dat_i[27]
port 296 nsew signal input
rlabel metal2 s 39144 74600 39200 75000 6 wb_dat_i[28]
port 297 nsew signal input
rlabel metal2 s 39760 74600 39816 75000 6 wb_dat_i[29]
port 298 nsew signal input
rlabel metal2 s 23128 74600 23184 75000 6 wb_dat_i[2]
port 299 nsew signal input
rlabel metal2 s 40376 74600 40432 75000 6 wb_dat_i[30]
port 300 nsew signal input
rlabel metal2 s 40992 74600 41048 75000 6 wb_dat_i[31]
port 301 nsew signal input
rlabel metal2 s 23744 74600 23800 75000 6 wb_dat_i[3]
port 302 nsew signal input
rlabel metal2 s 24360 74600 24416 75000 6 wb_dat_i[4]
port 303 nsew signal input
rlabel metal2 s 24976 74600 25032 75000 6 wb_dat_i[5]
port 304 nsew signal input
rlabel metal2 s 25592 74600 25648 75000 6 wb_dat_i[6]
port 305 nsew signal input
rlabel metal2 s 26208 74600 26264 75000 6 wb_dat_i[7]
port 306 nsew signal input
rlabel metal2 s 26824 74600 26880 75000 6 wb_dat_i[8]
port 307 nsew signal input
rlabel metal2 s 27440 74600 27496 75000 6 wb_dat_i[9]
port 308 nsew signal input
rlabel metal3 s 0 13104 400 13160 6 wb_dat_o[0]
port 309 nsew signal output
rlabel metal3 s 0 19264 400 19320 6 wb_dat_o[10]
port 310 nsew signal output
rlabel metal3 s 0 19880 400 19936 6 wb_dat_o[11]
port 311 nsew signal output
rlabel metal3 s 0 20496 400 20552 6 wb_dat_o[12]
port 312 nsew signal output
rlabel metal3 s 0 21112 400 21168 6 wb_dat_o[13]
port 313 nsew signal output
rlabel metal3 s 0 21728 400 21784 6 wb_dat_o[14]
port 314 nsew signal output
rlabel metal3 s 0 22344 400 22400 6 wb_dat_o[15]
port 315 nsew signal output
rlabel metal3 s 0 22960 400 23016 6 wb_dat_o[16]
port 316 nsew signal output
rlabel metal3 s 0 23576 400 23632 6 wb_dat_o[17]
port 317 nsew signal output
rlabel metal3 s 0 24192 400 24248 6 wb_dat_o[18]
port 318 nsew signal output
rlabel metal3 s 0 24808 400 24864 6 wb_dat_o[19]
port 319 nsew signal output
rlabel metal3 s 0 13720 400 13776 6 wb_dat_o[1]
port 320 nsew signal output
rlabel metal3 s 0 25424 400 25480 6 wb_dat_o[20]
port 321 nsew signal output
rlabel metal3 s 0 26040 400 26096 6 wb_dat_o[21]
port 322 nsew signal output
rlabel metal3 s 0 26656 400 26712 6 wb_dat_o[22]
port 323 nsew signal output
rlabel metal3 s 0 27272 400 27328 6 wb_dat_o[23]
port 324 nsew signal output
rlabel metal3 s 0 27888 400 27944 6 wb_dat_o[24]
port 325 nsew signal output
rlabel metal3 s 0 28504 400 28560 6 wb_dat_o[25]
port 326 nsew signal output
rlabel metal3 s 0 29120 400 29176 6 wb_dat_o[26]
port 327 nsew signal output
rlabel metal3 s 0 29736 400 29792 6 wb_dat_o[27]
port 328 nsew signal output
rlabel metal3 s 0 30352 400 30408 6 wb_dat_o[28]
port 329 nsew signal output
rlabel metal3 s 0 30968 400 31024 6 wb_dat_o[29]
port 330 nsew signal output
rlabel metal3 s 0 14336 400 14392 6 wb_dat_o[2]
port 331 nsew signal output
rlabel metal3 s 0 31584 400 31640 6 wb_dat_o[30]
port 332 nsew signal output
rlabel metal3 s 0 32200 400 32256 6 wb_dat_o[31]
port 333 nsew signal output
rlabel metal3 s 0 14952 400 15008 6 wb_dat_o[3]
port 334 nsew signal output
rlabel metal3 s 0 15568 400 15624 6 wb_dat_o[4]
port 335 nsew signal output
rlabel metal3 s 0 16184 400 16240 6 wb_dat_o[5]
port 336 nsew signal output
rlabel metal3 s 0 16800 400 16856 6 wb_dat_o[6]
port 337 nsew signal output
rlabel metal3 s 0 17416 400 17472 6 wb_dat_o[7]
port 338 nsew signal output
rlabel metal3 s 0 18032 400 18088 6 wb_dat_o[8]
port 339 nsew signal output
rlabel metal3 s 0 18648 400 18704 6 wb_dat_o[9]
port 340 nsew signal output
rlabel metal2 s 29232 0 29288 400 6 wb_rstn_i
port 341 nsew signal input
rlabel metal2 s 41608 74600 41664 75000 6 wb_sel_i[0]
port 342 nsew signal input
rlabel metal2 s 42224 74600 42280 75000 6 wb_sel_i[1]
port 343 nsew signal input
rlabel metal2 s 42840 74600 42896 75000 6 wb_sel_i[2]
port 344 nsew signal input
rlabel metal2 s 43456 74600 43512 75000 6 wb_sel_i[3]
port 345 nsew signal input
rlabel metal3 s 0 12488 400 12544 6 wb_stb_i
port 346 nsew signal input
rlabel metal2 s 44072 74600 44128 75000 6 wb_we_i
port 347 nsew signal input
<< properties >>
string FIXED_BBOX 0 0 47000 75000
string LEFclass BLOCK
string LEFview TRUE
string GDS_END 11723576
string GDS_FILE /home/hosni/GF180/caravel-gf180mcu/openlane/housekeeping/runs/RUN_2022.11.16_19.05.38/results/signoff/housekeeping.magic.gds
string GDS_START 566242
<< end >>

