VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO housekeeping
  CLASS BLOCK ;
  FOREIGN housekeeping ;
  ORIGIN 0.000 0.000 ;
  SIZE 470.000 BY 750.000 ;
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER Metal4 ;
        RECT 22.240 15.380 23.840 733.340 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 99.040 15.380 100.640 733.340 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 175.840 15.380 177.440 733.340 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 252.640 15.380 254.240 733.340 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 329.440 15.380 331.040 733.340 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 406.240 15.380 407.840 733.340 ;
    END
    PORT
      LAYER Metal5 ;
        RECT 6.420 31.290 463.420 32.890 ;
    END
    PORT
      LAYER Metal5 ;
        RECT 6.420 109.490 463.420 111.090 ;
    END
    PORT
      LAYER Metal5 ;
        RECT 6.420 187.690 463.420 189.290 ;
    END
    PORT
      LAYER Metal5 ;
        RECT 6.420 265.890 463.420 267.490 ;
    END
    PORT
      LAYER Metal5 ;
        RECT 6.420 344.090 463.420 345.690 ;
    END
    PORT
      LAYER Metal5 ;
        RECT 6.420 422.290 463.420 423.890 ;
    END
    PORT
      LAYER Metal5 ;
        RECT 6.420 500.490 463.420 502.090 ;
    END
    PORT
      LAYER Metal5 ;
        RECT 6.420 578.690 463.420 580.290 ;
    END
    PORT
      LAYER Metal5 ;
        RECT 6.420 656.890 463.420 658.490 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER Metal4 ;
        RECT 25.540 15.380 27.140 733.340 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 102.340 15.380 103.940 733.340 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 179.140 15.380 180.740 733.340 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 255.940 15.380 257.540 733.340 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 332.740 15.380 334.340 733.340 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 409.540 15.380 411.140 733.340 ;
    END
    PORT
      LAYER Metal5 ;
        RECT 6.420 70.390 463.420 71.990 ;
    END
    PORT
      LAYER Metal5 ;
        RECT 6.420 148.590 463.420 150.190 ;
    END
    PORT
      LAYER Metal5 ;
        RECT 6.420 226.790 463.420 228.390 ;
    END
    PORT
      LAYER Metal5 ;
        RECT 6.420 304.990 463.420 306.590 ;
    END
    PORT
      LAYER Metal5 ;
        RECT 6.420 383.190 463.420 384.790 ;
    END
    PORT
      LAYER Metal5 ;
        RECT 6.420 461.390 463.420 462.990 ;
    END
    PORT
      LAYER Metal5 ;
        RECT 6.420 539.590 463.420 541.190 ;
    END
    PORT
      LAYER Metal5 ;
        RECT 6.420 617.790 463.420 619.390 ;
    END
    PORT
      LAYER Metal5 ;
        RECT 6.420 695.990 463.420 697.590 ;
    END
  END VSS
  PIN debug_in
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 7.840 4.000 8.400 ;
    END
  END debug_in
  PIN debug_mode
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 14.000 4.000 14.560 ;
    END
  END debug_mode
  PIN debug_oeb
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 20.160 4.000 20.720 ;
    END
  END debug_oeb
  PIN debug_out
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 26.320 4.000 26.880 ;
    END
  END debug_out
  PIN irq[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 38.640 4.000 39.200 ;
    END
  END irq[0]
  PIN irq[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 44.800 4.000 45.360 ;
    END
  END irq[1]
  PIN irq[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 50.960 4.000 51.520 ;
    END
  END irq[2]
  PIN mask_rev_in[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 297.360 0.000 297.920 4.000 ;
    END
  END mask_rev_in[0]
  PIN mask_rev_in[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 347.760 0.000 348.320 4.000 ;
    END
  END mask_rev_in[10]
  PIN mask_rev_in[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 352.800 0.000 353.360 4.000 ;
    END
  END mask_rev_in[11]
  PIN mask_rev_in[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 357.840 0.000 358.400 4.000 ;
    END
  END mask_rev_in[12]
  PIN mask_rev_in[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 362.880 0.000 363.440 4.000 ;
    END
  END mask_rev_in[13]
  PIN mask_rev_in[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 367.920 0.000 368.480 4.000 ;
    END
  END mask_rev_in[14]
  PIN mask_rev_in[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 372.960 0.000 373.520 4.000 ;
    END
  END mask_rev_in[15]
  PIN mask_rev_in[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 378.000 0.000 378.560 4.000 ;
    END
  END mask_rev_in[16]
  PIN mask_rev_in[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 383.040 0.000 383.600 4.000 ;
    END
  END mask_rev_in[17]
  PIN mask_rev_in[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 388.080 0.000 388.640 4.000 ;
    END
  END mask_rev_in[18]
  PIN mask_rev_in[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 393.120 0.000 393.680 4.000 ;
    END
  END mask_rev_in[19]
  PIN mask_rev_in[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 302.400 0.000 302.960 4.000 ;
    END
  END mask_rev_in[1]
  PIN mask_rev_in[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 398.160 0.000 398.720 4.000 ;
    END
  END mask_rev_in[20]
  PIN mask_rev_in[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 403.200 0.000 403.760 4.000 ;
    END
  END mask_rev_in[21]
  PIN mask_rev_in[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 408.240 0.000 408.800 4.000 ;
    END
  END mask_rev_in[22]
  PIN mask_rev_in[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 413.280 0.000 413.840 4.000 ;
    END
  END mask_rev_in[23]
  PIN mask_rev_in[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 418.320 0.000 418.880 4.000 ;
    END
  END mask_rev_in[24]
  PIN mask_rev_in[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 423.360 0.000 423.920 4.000 ;
    END
  END mask_rev_in[25]
  PIN mask_rev_in[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 428.400 0.000 428.960 4.000 ;
    END
  END mask_rev_in[26]
  PIN mask_rev_in[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 433.440 0.000 434.000 4.000 ;
    END
  END mask_rev_in[27]
  PIN mask_rev_in[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 438.480 0.000 439.040 4.000 ;
    END
  END mask_rev_in[28]
  PIN mask_rev_in[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 443.520 0.000 444.080 4.000 ;
    END
  END mask_rev_in[29]
  PIN mask_rev_in[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 307.440 0.000 308.000 4.000 ;
    END
  END mask_rev_in[2]
  PIN mask_rev_in[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 448.560 0.000 449.120 4.000 ;
    END
  END mask_rev_in[30]
  PIN mask_rev_in[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 453.600 0.000 454.160 4.000 ;
    END
  END mask_rev_in[31]
  PIN mask_rev_in[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 312.480 0.000 313.040 4.000 ;
    END
  END mask_rev_in[3]
  PIN mask_rev_in[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 317.520 0.000 318.080 4.000 ;
    END
  END mask_rev_in[4]
  PIN mask_rev_in[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 322.560 0.000 323.120 4.000 ;
    END
  END mask_rev_in[5]
  PIN mask_rev_in[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 327.600 0.000 328.160 4.000 ;
    END
  END mask_rev_in[6]
  PIN mask_rev_in[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 332.640 0.000 333.200 4.000 ;
    END
  END mask_rev_in[7]
  PIN mask_rev_in[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 337.680 0.000 338.240 4.000 ;
    END
  END mask_rev_in[8]
  PIN mask_rev_in[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 342.720 0.000 343.280 4.000 ;
    END
  END mask_rev_in[9]
  PIN mgmt_gpio_in[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 466.000 72.240 470.000 72.800 ;
    END
  END mgmt_gpio_in[0]
  PIN mgmt_gpio_in[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 466.000 408.240 470.000 408.800 ;
    END
  END mgmt_gpio_in[10]
  PIN mgmt_gpio_in[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 466.000 441.840 470.000 442.400 ;
    END
  END mgmt_gpio_in[11]
  PIN mgmt_gpio_in[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 466.000 475.440 470.000 476.000 ;
    END
  END mgmt_gpio_in[12]
  PIN mgmt_gpio_in[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 466.000 509.040 470.000 509.600 ;
    END
  END mgmt_gpio_in[13]
  PIN mgmt_gpio_in[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 466.000 542.640 470.000 543.200 ;
    END
  END mgmt_gpio_in[14]
  PIN mgmt_gpio_in[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 466.000 576.240 470.000 576.800 ;
    END
  END mgmt_gpio_in[15]
  PIN mgmt_gpio_in[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 466.000 609.840 470.000 610.400 ;
    END
  END mgmt_gpio_in[16]
  PIN mgmt_gpio_in[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 466.000 643.440 470.000 644.000 ;
    END
  END mgmt_gpio_in[17]
  PIN mgmt_gpio_in[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 466.000 677.040 470.000 677.600 ;
    END
  END mgmt_gpio_in[18]
  PIN mgmt_gpio_in[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 466.000 710.640 470.000 711.200 ;
    END
  END mgmt_gpio_in[19]
  PIN mgmt_gpio_in[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 466.000 105.840 470.000 106.400 ;
    END
  END mgmt_gpio_in[1]
  PIN mgmt_gpio_in[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 414.400 4.000 414.960 ;
    END
  END mgmt_gpio_in[20]
  PIN mgmt_gpio_in[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 432.880 4.000 433.440 ;
    END
  END mgmt_gpio_in[21]
  PIN mgmt_gpio_in[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 451.360 4.000 451.920 ;
    END
  END mgmt_gpio_in[22]
  PIN mgmt_gpio_in[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 469.840 4.000 470.400 ;
    END
  END mgmt_gpio_in[23]
  PIN mgmt_gpio_in[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 488.320 4.000 488.880 ;
    END
  END mgmt_gpio_in[24]
  PIN mgmt_gpio_in[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 506.800 4.000 507.360 ;
    END
  END mgmt_gpio_in[25]
  PIN mgmt_gpio_in[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 525.280 4.000 525.840 ;
    END
  END mgmt_gpio_in[26]
  PIN mgmt_gpio_in[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 543.760 4.000 544.320 ;
    END
  END mgmt_gpio_in[27]
  PIN mgmt_gpio_in[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 562.240 4.000 562.800 ;
    END
  END mgmt_gpio_in[28]
  PIN mgmt_gpio_in[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 580.720 4.000 581.280 ;
    END
  END mgmt_gpio_in[29]
  PIN mgmt_gpio_in[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 466.000 139.440 470.000 140.000 ;
    END
  END mgmt_gpio_in[2]
  PIN mgmt_gpio_in[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 599.200 4.000 599.760 ;
    END
  END mgmt_gpio_in[30]
  PIN mgmt_gpio_in[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 617.680 4.000 618.240 ;
    END
  END mgmt_gpio_in[31]
  PIN mgmt_gpio_in[32]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 636.160 4.000 636.720 ;
    END
  END mgmt_gpio_in[32]
  PIN mgmt_gpio_in[33]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 654.640 4.000 655.200 ;
    END
  END mgmt_gpio_in[33]
  PIN mgmt_gpio_in[34]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 673.120 4.000 673.680 ;
    END
  END mgmt_gpio_in[34]
  PIN mgmt_gpio_in[35]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 691.600 4.000 692.160 ;
    END
  END mgmt_gpio_in[35]
  PIN mgmt_gpio_in[36]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 710.080 4.000 710.640 ;
    END
  END mgmt_gpio_in[36]
  PIN mgmt_gpio_in[37]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 728.560 4.000 729.120 ;
    END
  END mgmt_gpio_in[37]
  PIN mgmt_gpio_in[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 466.000 173.040 470.000 173.600 ;
    END
  END mgmt_gpio_in[3]
  PIN mgmt_gpio_in[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 466.000 206.640 470.000 207.200 ;
    END
  END mgmt_gpio_in[4]
  PIN mgmt_gpio_in[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 466.000 240.240 470.000 240.800 ;
    END
  END mgmt_gpio_in[5]
  PIN mgmt_gpio_in[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 466.000 273.840 470.000 274.400 ;
    END
  END mgmt_gpio_in[6]
  PIN mgmt_gpio_in[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 466.000 307.440 470.000 308.000 ;
    END
  END mgmt_gpio_in[7]
  PIN mgmt_gpio_in[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 466.000 341.040 470.000 341.600 ;
    END
  END mgmt_gpio_in[8]
  PIN mgmt_gpio_in[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 466.000 374.640 470.000 375.200 ;
    END
  END mgmt_gpio_in[9]
  PIN mgmt_gpio_oeb[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 466.000 83.440 470.000 84.000 ;
    END
  END mgmt_gpio_oeb[0]
  PIN mgmt_gpio_oeb[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 466.000 419.440 470.000 420.000 ;
    END
  END mgmt_gpio_oeb[10]
  PIN mgmt_gpio_oeb[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 466.000 453.040 470.000 453.600 ;
    END
  END mgmt_gpio_oeb[11]
  PIN mgmt_gpio_oeb[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 466.000 486.640 470.000 487.200 ;
    END
  END mgmt_gpio_oeb[12]
  PIN mgmt_gpio_oeb[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 466.000 520.240 470.000 520.800 ;
    END
  END mgmt_gpio_oeb[13]
  PIN mgmt_gpio_oeb[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 466.000 553.840 470.000 554.400 ;
    END
  END mgmt_gpio_oeb[14]
  PIN mgmt_gpio_oeb[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 466.000 587.440 470.000 588.000 ;
    END
  END mgmt_gpio_oeb[15]
  PIN mgmt_gpio_oeb[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 466.000 621.040 470.000 621.600 ;
    END
  END mgmt_gpio_oeb[16]
  PIN mgmt_gpio_oeb[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 466.000 654.640 470.000 655.200 ;
    END
  END mgmt_gpio_oeb[17]
  PIN mgmt_gpio_oeb[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 466.000 688.240 470.000 688.800 ;
    END
  END mgmt_gpio_oeb[18]
  PIN mgmt_gpio_oeb[19]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 466.000 721.840 470.000 722.400 ;
    END
  END mgmt_gpio_oeb[19]
  PIN mgmt_gpio_oeb[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 466.000 117.040 470.000 117.600 ;
    END
  END mgmt_gpio_oeb[1]
  PIN mgmt_gpio_oeb[20]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 420.560 4.000 421.120 ;
    END
  END mgmt_gpio_oeb[20]
  PIN mgmt_gpio_oeb[21]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 439.040 4.000 439.600 ;
    END
  END mgmt_gpio_oeb[21]
  PIN mgmt_gpio_oeb[22]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 457.520 4.000 458.080 ;
    END
  END mgmt_gpio_oeb[22]
  PIN mgmt_gpio_oeb[23]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 476.000 4.000 476.560 ;
    END
  END mgmt_gpio_oeb[23]
  PIN mgmt_gpio_oeb[24]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 494.480 4.000 495.040 ;
    END
  END mgmt_gpio_oeb[24]
  PIN mgmt_gpio_oeb[25]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 512.960 4.000 513.520 ;
    END
  END mgmt_gpio_oeb[25]
  PIN mgmt_gpio_oeb[26]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 531.440 4.000 532.000 ;
    END
  END mgmt_gpio_oeb[26]
  PIN mgmt_gpio_oeb[27]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 549.920 4.000 550.480 ;
    END
  END mgmt_gpio_oeb[27]
  PIN mgmt_gpio_oeb[28]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 568.400 4.000 568.960 ;
    END
  END mgmt_gpio_oeb[28]
  PIN mgmt_gpio_oeb[29]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 586.880 4.000 587.440 ;
    END
  END mgmt_gpio_oeb[29]
  PIN mgmt_gpio_oeb[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 466.000 150.640 470.000 151.200 ;
    END
  END mgmt_gpio_oeb[2]
  PIN mgmt_gpio_oeb[30]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 605.360 4.000 605.920 ;
    END
  END mgmt_gpio_oeb[30]
  PIN mgmt_gpio_oeb[31]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 623.840 4.000 624.400 ;
    END
  END mgmt_gpio_oeb[31]
  PIN mgmt_gpio_oeb[32]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 642.320 4.000 642.880 ;
    END
  END mgmt_gpio_oeb[32]
  PIN mgmt_gpio_oeb[33]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 660.800 4.000 661.360 ;
    END
  END mgmt_gpio_oeb[33]
  PIN mgmt_gpio_oeb[34]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 679.280 4.000 679.840 ;
    END
  END mgmt_gpio_oeb[34]
  PIN mgmt_gpio_oeb[35]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 697.760 4.000 698.320 ;
    END
  END mgmt_gpio_oeb[35]
  PIN mgmt_gpio_oeb[36]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 716.240 4.000 716.800 ;
    END
  END mgmt_gpio_oeb[36]
  PIN mgmt_gpio_oeb[37]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 734.720 4.000 735.280 ;
    END
  END mgmt_gpio_oeb[37]
  PIN mgmt_gpio_oeb[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 466.000 184.240 470.000 184.800 ;
    END
  END mgmt_gpio_oeb[3]
  PIN mgmt_gpio_oeb[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 466.000 217.840 470.000 218.400 ;
    END
  END mgmt_gpio_oeb[4]
  PIN mgmt_gpio_oeb[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 466.000 251.440 470.000 252.000 ;
    END
  END mgmt_gpio_oeb[5]
  PIN mgmt_gpio_oeb[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 466.000 285.040 470.000 285.600 ;
    END
  END mgmt_gpio_oeb[6]
  PIN mgmt_gpio_oeb[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 466.000 318.640 470.000 319.200 ;
    END
  END mgmt_gpio_oeb[7]
  PIN mgmt_gpio_oeb[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 466.000 352.240 470.000 352.800 ;
    END
  END mgmt_gpio_oeb[8]
  PIN mgmt_gpio_oeb[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 466.000 385.840 470.000 386.400 ;
    END
  END mgmt_gpio_oeb[9]
  PIN mgmt_gpio_out[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 466.000 94.640 470.000 95.200 ;
    END
  END mgmt_gpio_out[0]
  PIN mgmt_gpio_out[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 466.000 430.640 470.000 431.200 ;
    END
  END mgmt_gpio_out[10]
  PIN mgmt_gpio_out[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 466.000 464.240 470.000 464.800 ;
    END
  END mgmt_gpio_out[11]
  PIN mgmt_gpio_out[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 466.000 497.840 470.000 498.400 ;
    END
  END mgmt_gpio_out[12]
  PIN mgmt_gpio_out[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 466.000 531.440 470.000 532.000 ;
    END
  END mgmt_gpio_out[13]
  PIN mgmt_gpio_out[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 466.000 565.040 470.000 565.600 ;
    END
  END mgmt_gpio_out[14]
  PIN mgmt_gpio_out[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 466.000 598.640 470.000 599.200 ;
    END
  END mgmt_gpio_out[15]
  PIN mgmt_gpio_out[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 466.000 632.240 470.000 632.800 ;
    END
  END mgmt_gpio_out[16]
  PIN mgmt_gpio_out[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 466.000 665.840 470.000 666.400 ;
    END
  END mgmt_gpio_out[17]
  PIN mgmt_gpio_out[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 466.000 699.440 470.000 700.000 ;
    END
  END mgmt_gpio_out[18]
  PIN mgmt_gpio_out[19]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 466.000 733.040 470.000 733.600 ;
    END
  END mgmt_gpio_out[19]
  PIN mgmt_gpio_out[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 466.000 128.240 470.000 128.800 ;
    END
  END mgmt_gpio_out[1]
  PIN mgmt_gpio_out[20]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 426.720 4.000 427.280 ;
    END
  END mgmt_gpio_out[20]
  PIN mgmt_gpio_out[21]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 445.200 4.000 445.760 ;
    END
  END mgmt_gpio_out[21]
  PIN mgmt_gpio_out[22]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 463.680 4.000 464.240 ;
    END
  END mgmt_gpio_out[22]
  PIN mgmt_gpio_out[23]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 482.160 4.000 482.720 ;
    END
  END mgmt_gpio_out[23]
  PIN mgmt_gpio_out[24]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 500.640 4.000 501.200 ;
    END
  END mgmt_gpio_out[24]
  PIN mgmt_gpio_out[25]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 519.120 4.000 519.680 ;
    END
  END mgmt_gpio_out[25]
  PIN mgmt_gpio_out[26]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 537.600 4.000 538.160 ;
    END
  END mgmt_gpio_out[26]
  PIN mgmt_gpio_out[27]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 556.080 4.000 556.640 ;
    END
  END mgmt_gpio_out[27]
  PIN mgmt_gpio_out[28]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 574.560 4.000 575.120 ;
    END
  END mgmt_gpio_out[28]
  PIN mgmt_gpio_out[29]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 593.040 4.000 593.600 ;
    END
  END mgmt_gpio_out[29]
  PIN mgmt_gpio_out[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 466.000 161.840 470.000 162.400 ;
    END
  END mgmt_gpio_out[2]
  PIN mgmt_gpio_out[30]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 611.520 4.000 612.080 ;
    END
  END mgmt_gpio_out[30]
  PIN mgmt_gpio_out[31]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 630.000 4.000 630.560 ;
    END
  END mgmt_gpio_out[31]
  PIN mgmt_gpio_out[32]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 648.480 4.000 649.040 ;
    END
  END mgmt_gpio_out[32]
  PIN mgmt_gpio_out[33]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 666.960 4.000 667.520 ;
    END
  END mgmt_gpio_out[33]
  PIN mgmt_gpio_out[34]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 685.440 4.000 686.000 ;
    END
  END mgmt_gpio_out[34]
  PIN mgmt_gpio_out[35]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 703.920 4.000 704.480 ;
    END
  END mgmt_gpio_out[35]
  PIN mgmt_gpio_out[36]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 722.400 4.000 722.960 ;
    END
  END mgmt_gpio_out[36]
  PIN mgmt_gpio_out[37]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 740.880 4.000 741.440 ;
    END
  END mgmt_gpio_out[37]
  PIN mgmt_gpio_out[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 466.000 195.440 470.000 196.000 ;
    END
  END mgmt_gpio_out[3]
  PIN mgmt_gpio_out[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 466.000 229.040 470.000 229.600 ;
    END
  END mgmt_gpio_out[4]
  PIN mgmt_gpio_out[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 466.000 262.640 470.000 263.200 ;
    END
  END mgmt_gpio_out[5]
  PIN mgmt_gpio_out[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 466.000 296.240 470.000 296.800 ;
    END
  END mgmt_gpio_out[6]
  PIN mgmt_gpio_out[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 466.000 329.840 470.000 330.400 ;
    END
  END mgmt_gpio_out[7]
  PIN mgmt_gpio_out[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 466.000 363.440 470.000 364.000 ;
    END
  END mgmt_gpio_out[8]
  PIN mgmt_gpio_out[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 466.000 397.040 470.000 397.600 ;
    END
  END mgmt_gpio_out[9]
  PIN pad_flash_clk
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 15.120 0.000 15.680 4.000 ;
    END
  END pad_flash_clk
  PIN pad_flash_clk_oe
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 20.160 0.000 20.720 4.000 ;
    END
  END pad_flash_clk_oe
  PIN pad_flash_csb
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 25.200 0.000 25.760 4.000 ;
    END
  END pad_flash_csb
  PIN pad_flash_csb_oe
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 30.240 0.000 30.800 4.000 ;
    END
  END pad_flash_csb_oe
  PIN pad_flash_io0_di
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 35.280 0.000 35.840 4.000 ;
    END
  END pad_flash_io0_di
  PIN pad_flash_io0_do
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 40.320 0.000 40.880 4.000 ;
    END
  END pad_flash_io0_do
  PIN pad_flash_io0_ie
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 45.360 0.000 45.920 4.000 ;
    END
  END pad_flash_io0_ie
  PIN pad_flash_io0_oe
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 50.400 0.000 50.960 4.000 ;
    END
  END pad_flash_io0_oe
  PIN pad_flash_io1_di
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 55.440 0.000 56.000 4.000 ;
    END
  END pad_flash_io1_di
  PIN pad_flash_io1_do
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 60.480 0.000 61.040 4.000 ;
    END
  END pad_flash_io1_do
  PIN pad_flash_io1_ie
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 65.520 0.000 66.080 4.000 ;
    END
  END pad_flash_io1_ie
  PIN pad_flash_io1_oe
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 70.560 0.000 71.120 4.000 ;
    END
  END pad_flash_io1_oe
  PIN pll90_sel[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 136.080 0.000 136.640 4.000 ;
    END
  END pll90_sel[0]
  PIN pll90_sel[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 141.120 0.000 141.680 4.000 ;
    END
  END pll90_sel[1]
  PIN pll90_sel[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 146.160 0.000 146.720 4.000 ;
    END
  END pll90_sel[2]
  PIN pll_bypass
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 282.240 0.000 282.800 4.000 ;
    END
  END pll_bypass
  PIN pll_dco_ena
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 90.720 0.000 91.280 4.000 ;
    END
  END pll_dco_ena
  PIN pll_div[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 95.760 0.000 96.320 4.000 ;
    END
  END pll_div[0]
  PIN pll_div[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 100.800 0.000 101.360 4.000 ;
    END
  END pll_div[1]
  PIN pll_div[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 105.840 0.000 106.400 4.000 ;
    END
  END pll_div[2]
  PIN pll_div[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 110.880 0.000 111.440 4.000 ;
    END
  END pll_div[3]
  PIN pll_div[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 115.920 0.000 116.480 4.000 ;
    END
  END pll_div[4]
  PIN pll_ena
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 85.680 0.000 86.240 4.000 ;
    END
  END pll_ena
  PIN pll_sel[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 120.960 0.000 121.520 4.000 ;
    END
  END pll_sel[0]
  PIN pll_sel[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 126.000 0.000 126.560 4.000 ;
    END
  END pll_sel[1]
  PIN pll_sel[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 131.040 0.000 131.600 4.000 ;
    END
  END pll_sel[2]
  PIN pll_trim[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 151.200 0.000 151.760 4.000 ;
    END
  END pll_trim[0]
  PIN pll_trim[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 201.600 0.000 202.160 4.000 ;
    END
  END pll_trim[10]
  PIN pll_trim[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 206.640 0.000 207.200 4.000 ;
    END
  END pll_trim[11]
  PIN pll_trim[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 211.680 0.000 212.240 4.000 ;
    END
  END pll_trim[12]
  PIN pll_trim[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 216.720 0.000 217.280 4.000 ;
    END
  END pll_trim[13]
  PIN pll_trim[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 221.760 0.000 222.320 4.000 ;
    END
  END pll_trim[14]
  PIN pll_trim[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 226.800 0.000 227.360 4.000 ;
    END
  END pll_trim[15]
  PIN pll_trim[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 231.840 0.000 232.400 4.000 ;
    END
  END pll_trim[16]
  PIN pll_trim[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 236.880 0.000 237.440 4.000 ;
    END
  END pll_trim[17]
  PIN pll_trim[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 241.920 0.000 242.480 4.000 ;
    END
  END pll_trim[18]
  PIN pll_trim[19]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 246.960 0.000 247.520 4.000 ;
    END
  END pll_trim[19]
  PIN pll_trim[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 156.240 0.000 156.800 4.000 ;
    END
  END pll_trim[1]
  PIN pll_trim[20]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 252.000 0.000 252.560 4.000 ;
    END
  END pll_trim[20]
  PIN pll_trim[21]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 257.040 0.000 257.600 4.000 ;
    END
  END pll_trim[21]
  PIN pll_trim[22]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 262.080 0.000 262.640 4.000 ;
    END
  END pll_trim[22]
  PIN pll_trim[23]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 267.120 0.000 267.680 4.000 ;
    END
  END pll_trim[23]
  PIN pll_trim[24]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 272.160 0.000 272.720 4.000 ;
    END
  END pll_trim[24]
  PIN pll_trim[25]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 277.200 0.000 277.760 4.000 ;
    END
  END pll_trim[25]
  PIN pll_trim[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 161.280 0.000 161.840 4.000 ;
    END
  END pll_trim[2]
  PIN pll_trim[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 166.320 0.000 166.880 4.000 ;
    END
  END pll_trim[3]
  PIN pll_trim[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 171.360 0.000 171.920 4.000 ;
    END
  END pll_trim[4]
  PIN pll_trim[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 176.400 0.000 176.960 4.000 ;
    END
  END pll_trim[5]
  PIN pll_trim[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 181.440 0.000 182.000 4.000 ;
    END
  END pll_trim[6]
  PIN pll_trim[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 186.480 0.000 187.040 4.000 ;
    END
  END pll_trim[7]
  PIN pll_trim[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 191.520 0.000 192.080 4.000 ;
    END
  END pll_trim[8]
  PIN pll_trim[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 196.560 0.000 197.120 4.000 ;
    END
  END pll_trim[9]
  PIN porb
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 75.600 0.000 76.160 4.000 ;
    END
  END porb
  PIN pwr_ctrl_out
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 458.640 0.000 459.200 4.000 ;
    END
  END pwr_ctrl_out
  PIN qspi_enabled
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 100.240 4.000 100.800 ;
    END
  END qspi_enabled
  PIN reset
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 80.640 0.000 81.200 4.000 ;
    END
  END reset
  PIN ser_rx
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 94.080 4.000 94.640 ;
    END
  END ser_rx
  PIN ser_tx
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 87.920 4.000 88.480 ;
    END
  END ser_tx
  PIN serial_clock
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 466.000 16.240 470.000 16.800 ;
    END
  END serial_clock
  PIN serial_data_1
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 466.000 49.840 470.000 50.400 ;
    END
  END serial_data_1
  PIN serial_data_2
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 466.000 61.040 470.000 61.600 ;
    END
  END serial_data_2
  PIN serial_load
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 466.000 38.640 470.000 39.200 ;
    END
  END serial_load
  PIN serial_resetn
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 466.000 27.440 470.000 28.000 ;
    END
  END serial_resetn
  PIN spi_csb
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 75.600 4.000 76.160 ;
    END
  END spi_csb
  PIN spi_enabled
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 112.560 4.000 113.120 ;
    END
  END spi_enabled
  PIN spi_sck
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 69.440 4.000 70.000 ;
    END
  END spi_sck
  PIN spi_sdi
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 81.760 4.000 82.320 ;
    END
  END spi_sdi
  PIN spi_sdo
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 63.280 4.000 63.840 ;
    END
  END spi_sdo
  PIN spi_sdoenb
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 57.120 4.000 57.680 ;
    END
  END spi_sdoenb
  PIN spimemio_flash_clk
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 328.160 4.000 328.720 ;
    END
  END spimemio_flash_clk
  PIN spimemio_flash_csb
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 334.320 4.000 334.880 ;
    END
  END spimemio_flash_csb
  PIN spimemio_flash_io0_di
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 340.480 4.000 341.040 ;
    END
  END spimemio_flash_io0_di
  PIN spimemio_flash_io0_do
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 346.640 4.000 347.200 ;
    END
  END spimemio_flash_io0_do
  PIN spimemio_flash_io0_oeb
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 352.800 4.000 353.360 ;
    END
  END spimemio_flash_io0_oeb
  PIN spimemio_flash_io1_di
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 358.960 4.000 359.520 ;
    END
  END spimemio_flash_io1_di
  PIN spimemio_flash_io1_do
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 365.120 4.000 365.680 ;
    END
  END spimemio_flash_io1_do
  PIN spimemio_flash_io1_oeb
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 371.280 4.000 371.840 ;
    END
  END spimemio_flash_io1_oeb
  PIN spimemio_flash_io2_di
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 377.440 4.000 378.000 ;
    END
  END spimemio_flash_io2_di
  PIN spimemio_flash_io2_do
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 383.600 4.000 384.160 ;
    END
  END spimemio_flash_io2_do
  PIN spimemio_flash_io2_oeb
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 389.760 4.000 390.320 ;
    END
  END spimemio_flash_io2_oeb
  PIN spimemio_flash_io3_di
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 395.920 4.000 396.480 ;
    END
  END spimemio_flash_io3_di
  PIN spimemio_flash_io3_do
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 402.080 4.000 402.640 ;
    END
  END spimemio_flash_io3_do
  PIN spimemio_flash_io3_oeb
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 408.240 4.000 408.800 ;
    END
  END spimemio_flash_io3_oeb
  PIN trap
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 32.480 4.000 33.040 ;
    END
  END trap
  PIN uart_enabled
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 106.400 4.000 106.960 ;
    END
  END uart_enabled
  PIN user_clock
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 10.080 0.000 10.640 4.000 ;
    END
  END user_clock
  PIN wb_ack_o
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 118.720 4.000 119.280 ;
    END
  END wb_ack_o
  PIN wb_adr_i[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 21.840 746.000 22.400 750.000 ;
    END
  END wb_adr_i[0]
  PIN wb_adr_i[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 83.440 746.000 84.000 750.000 ;
    END
  END wb_adr_i[10]
  PIN wb_adr_i[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 89.600 746.000 90.160 750.000 ;
    END
  END wb_adr_i[11]
  PIN wb_adr_i[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 95.760 746.000 96.320 750.000 ;
    END
  END wb_adr_i[12]
  PIN wb_adr_i[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 101.920 746.000 102.480 750.000 ;
    END
  END wb_adr_i[13]
  PIN wb_adr_i[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 108.080 746.000 108.640 750.000 ;
    END
  END wb_adr_i[14]
  PIN wb_adr_i[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 114.240 746.000 114.800 750.000 ;
    END
  END wb_adr_i[15]
  PIN wb_adr_i[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 120.400 746.000 120.960 750.000 ;
    END
  END wb_adr_i[16]
  PIN wb_adr_i[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 126.560 746.000 127.120 750.000 ;
    END
  END wb_adr_i[17]
  PIN wb_adr_i[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 132.720 746.000 133.280 750.000 ;
    END
  END wb_adr_i[18]
  PIN wb_adr_i[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 138.880 746.000 139.440 750.000 ;
    END
  END wb_adr_i[19]
  PIN wb_adr_i[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 28.000 746.000 28.560 750.000 ;
    END
  END wb_adr_i[1]
  PIN wb_adr_i[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 145.040 746.000 145.600 750.000 ;
    END
  END wb_adr_i[20]
  PIN wb_adr_i[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 151.200 746.000 151.760 750.000 ;
    END
  END wb_adr_i[21]
  PIN wb_adr_i[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 157.360 746.000 157.920 750.000 ;
    END
  END wb_adr_i[22]
  PIN wb_adr_i[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 163.520 746.000 164.080 750.000 ;
    END
  END wb_adr_i[23]
  PIN wb_adr_i[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 169.680 746.000 170.240 750.000 ;
    END
  END wb_adr_i[24]
  PIN wb_adr_i[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 175.840 746.000 176.400 750.000 ;
    END
  END wb_adr_i[25]
  PIN wb_adr_i[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 182.000 746.000 182.560 750.000 ;
    END
  END wb_adr_i[26]
  PIN wb_adr_i[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 188.160 746.000 188.720 750.000 ;
    END
  END wb_adr_i[27]
  PIN wb_adr_i[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 194.320 746.000 194.880 750.000 ;
    END
  END wb_adr_i[28]
  PIN wb_adr_i[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 200.480 746.000 201.040 750.000 ;
    END
  END wb_adr_i[29]
  PIN wb_adr_i[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 34.160 746.000 34.720 750.000 ;
    END
  END wb_adr_i[2]
  PIN wb_adr_i[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 206.640 746.000 207.200 750.000 ;
    END
  END wb_adr_i[30]
  PIN wb_adr_i[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 212.800 746.000 213.360 750.000 ;
    END
  END wb_adr_i[31]
  PIN wb_adr_i[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 40.320 746.000 40.880 750.000 ;
    END
  END wb_adr_i[3]
  PIN wb_adr_i[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 46.480 746.000 47.040 750.000 ;
    END
  END wb_adr_i[4]
  PIN wb_adr_i[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 52.640 746.000 53.200 750.000 ;
    END
  END wb_adr_i[5]
  PIN wb_adr_i[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 58.800 746.000 59.360 750.000 ;
    END
  END wb_adr_i[6]
  PIN wb_adr_i[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 64.960 746.000 65.520 750.000 ;
    END
  END wb_adr_i[7]
  PIN wb_adr_i[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 71.120 746.000 71.680 750.000 ;
    END
  END wb_adr_i[8]
  PIN wb_adr_i[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 77.280 746.000 77.840 750.000 ;
    END
  END wb_adr_i[9]
  PIN wb_clk_i
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 287.280 0.000 287.840 4.000 ;
    END
  END wb_clk_i
  PIN wb_cyc_i
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 446.880 746.000 447.440 750.000 ;
    END
  END wb_cyc_i
  PIN wb_dat_i[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 218.960 746.000 219.520 750.000 ;
    END
  END wb_dat_i[0]
  PIN wb_dat_i[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 280.560 746.000 281.120 750.000 ;
    END
  END wb_dat_i[10]
  PIN wb_dat_i[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 286.720 746.000 287.280 750.000 ;
    END
  END wb_dat_i[11]
  PIN wb_dat_i[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 292.880 746.000 293.440 750.000 ;
    END
  END wb_dat_i[12]
  PIN wb_dat_i[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 299.040 746.000 299.600 750.000 ;
    END
  END wb_dat_i[13]
  PIN wb_dat_i[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 305.200 746.000 305.760 750.000 ;
    END
  END wb_dat_i[14]
  PIN wb_dat_i[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 311.360 746.000 311.920 750.000 ;
    END
  END wb_dat_i[15]
  PIN wb_dat_i[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 317.520 746.000 318.080 750.000 ;
    END
  END wb_dat_i[16]
  PIN wb_dat_i[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 323.680 746.000 324.240 750.000 ;
    END
  END wb_dat_i[17]
  PIN wb_dat_i[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 329.840 746.000 330.400 750.000 ;
    END
  END wb_dat_i[18]
  PIN wb_dat_i[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 336.000 746.000 336.560 750.000 ;
    END
  END wb_dat_i[19]
  PIN wb_dat_i[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 225.120 746.000 225.680 750.000 ;
    END
  END wb_dat_i[1]
  PIN wb_dat_i[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 342.160 746.000 342.720 750.000 ;
    END
  END wb_dat_i[20]
  PIN wb_dat_i[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 348.320 746.000 348.880 750.000 ;
    END
  END wb_dat_i[21]
  PIN wb_dat_i[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 354.480 746.000 355.040 750.000 ;
    END
  END wb_dat_i[22]
  PIN wb_dat_i[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 360.640 746.000 361.200 750.000 ;
    END
  END wb_dat_i[23]
  PIN wb_dat_i[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 366.800 746.000 367.360 750.000 ;
    END
  END wb_dat_i[24]
  PIN wb_dat_i[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 372.960 746.000 373.520 750.000 ;
    END
  END wb_dat_i[25]
  PIN wb_dat_i[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 379.120 746.000 379.680 750.000 ;
    END
  END wb_dat_i[26]
  PIN wb_dat_i[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 385.280 746.000 385.840 750.000 ;
    END
  END wb_dat_i[27]
  PIN wb_dat_i[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 391.440 746.000 392.000 750.000 ;
    END
  END wb_dat_i[28]
  PIN wb_dat_i[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 397.600 746.000 398.160 750.000 ;
    END
  END wb_dat_i[29]
  PIN wb_dat_i[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 231.280 746.000 231.840 750.000 ;
    END
  END wb_dat_i[2]
  PIN wb_dat_i[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 403.760 746.000 404.320 750.000 ;
    END
  END wb_dat_i[30]
  PIN wb_dat_i[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 409.920 746.000 410.480 750.000 ;
    END
  END wb_dat_i[31]
  PIN wb_dat_i[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 237.440 746.000 238.000 750.000 ;
    END
  END wb_dat_i[3]
  PIN wb_dat_i[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 243.600 746.000 244.160 750.000 ;
    END
  END wb_dat_i[4]
  PIN wb_dat_i[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 249.760 746.000 250.320 750.000 ;
    END
  END wb_dat_i[5]
  PIN wb_dat_i[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 255.920 746.000 256.480 750.000 ;
    END
  END wb_dat_i[6]
  PIN wb_dat_i[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 262.080 746.000 262.640 750.000 ;
    END
  END wb_dat_i[7]
  PIN wb_dat_i[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 268.240 746.000 268.800 750.000 ;
    END
  END wb_dat_i[8]
  PIN wb_dat_i[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 274.400 746.000 274.960 750.000 ;
    END
  END wb_dat_i[9]
  PIN wb_dat_o[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 131.040 4.000 131.600 ;
    END
  END wb_dat_o[0]
  PIN wb_dat_o[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 192.640 4.000 193.200 ;
    END
  END wb_dat_o[10]
  PIN wb_dat_o[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 198.800 4.000 199.360 ;
    END
  END wb_dat_o[11]
  PIN wb_dat_o[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 204.960 4.000 205.520 ;
    END
  END wb_dat_o[12]
  PIN wb_dat_o[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 211.120 4.000 211.680 ;
    END
  END wb_dat_o[13]
  PIN wb_dat_o[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 217.280 4.000 217.840 ;
    END
  END wb_dat_o[14]
  PIN wb_dat_o[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 223.440 4.000 224.000 ;
    END
  END wb_dat_o[15]
  PIN wb_dat_o[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 229.600 4.000 230.160 ;
    END
  END wb_dat_o[16]
  PIN wb_dat_o[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 235.760 4.000 236.320 ;
    END
  END wb_dat_o[17]
  PIN wb_dat_o[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 241.920 4.000 242.480 ;
    END
  END wb_dat_o[18]
  PIN wb_dat_o[19]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 248.080 4.000 248.640 ;
    END
  END wb_dat_o[19]
  PIN wb_dat_o[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 137.200 4.000 137.760 ;
    END
  END wb_dat_o[1]
  PIN wb_dat_o[20]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 254.240 4.000 254.800 ;
    END
  END wb_dat_o[20]
  PIN wb_dat_o[21]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 260.400 4.000 260.960 ;
    END
  END wb_dat_o[21]
  PIN wb_dat_o[22]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 266.560 4.000 267.120 ;
    END
  END wb_dat_o[22]
  PIN wb_dat_o[23]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 272.720 4.000 273.280 ;
    END
  END wb_dat_o[23]
  PIN wb_dat_o[24]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 278.880 4.000 279.440 ;
    END
  END wb_dat_o[24]
  PIN wb_dat_o[25]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 285.040 4.000 285.600 ;
    END
  END wb_dat_o[25]
  PIN wb_dat_o[26]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 291.200 4.000 291.760 ;
    END
  END wb_dat_o[26]
  PIN wb_dat_o[27]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 297.360 4.000 297.920 ;
    END
  END wb_dat_o[27]
  PIN wb_dat_o[28]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 303.520 4.000 304.080 ;
    END
  END wb_dat_o[28]
  PIN wb_dat_o[29]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 309.680 4.000 310.240 ;
    END
  END wb_dat_o[29]
  PIN wb_dat_o[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 143.360 4.000 143.920 ;
    END
  END wb_dat_o[2]
  PIN wb_dat_o[30]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 315.840 4.000 316.400 ;
    END
  END wb_dat_o[30]
  PIN wb_dat_o[31]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 322.000 4.000 322.560 ;
    END
  END wb_dat_o[31]
  PIN wb_dat_o[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 149.520 4.000 150.080 ;
    END
  END wb_dat_o[3]
  PIN wb_dat_o[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 155.680 4.000 156.240 ;
    END
  END wb_dat_o[4]
  PIN wb_dat_o[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 161.840 4.000 162.400 ;
    END
  END wb_dat_o[5]
  PIN wb_dat_o[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 168.000 4.000 168.560 ;
    END
  END wb_dat_o[6]
  PIN wb_dat_o[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 174.160 4.000 174.720 ;
    END
  END wb_dat_o[7]
  PIN wb_dat_o[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 180.320 4.000 180.880 ;
    END
  END wb_dat_o[8]
  PIN wb_dat_o[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 186.480 4.000 187.040 ;
    END
  END wb_dat_o[9]
  PIN wb_rstn_i
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 292.320 0.000 292.880 4.000 ;
    END
  END wb_rstn_i
  PIN wb_sel_i[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 416.080 746.000 416.640 750.000 ;
    END
  END wb_sel_i[0]
  PIN wb_sel_i[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 422.240 746.000 422.800 750.000 ;
    END
  END wb_sel_i[1]
  PIN wb_sel_i[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 428.400 746.000 428.960 750.000 ;
    END
  END wb_sel_i[2]
  PIN wb_sel_i[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 434.560 746.000 435.120 750.000 ;
    END
  END wb_sel_i[3]
  PIN wb_stb_i
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 124.880 4.000 125.440 ;
    END
  END wb_stb_i
  PIN wb_we_i
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 440.720 746.000 441.280 750.000 ;
    END
  END wb_we_i
  OBS
      LAYER Metal1 ;
        RECT 6.720 15.380 469.750 734.010 ;
      LAYER Metal2 ;
        RECT 7.420 745.700 21.540 749.750 ;
        RECT 22.700 745.700 27.700 749.750 ;
        RECT 28.860 745.700 33.860 749.750 ;
        RECT 35.020 745.700 40.020 749.750 ;
        RECT 41.180 745.700 46.180 749.750 ;
        RECT 47.340 745.700 52.340 749.750 ;
        RECT 53.500 745.700 58.500 749.750 ;
        RECT 59.660 745.700 64.660 749.750 ;
        RECT 65.820 745.700 70.820 749.750 ;
        RECT 71.980 745.700 76.980 749.750 ;
        RECT 78.140 745.700 83.140 749.750 ;
        RECT 84.300 745.700 89.300 749.750 ;
        RECT 90.460 745.700 95.460 749.750 ;
        RECT 96.620 745.700 101.620 749.750 ;
        RECT 102.780 745.700 107.780 749.750 ;
        RECT 108.940 745.700 113.940 749.750 ;
        RECT 115.100 745.700 120.100 749.750 ;
        RECT 121.260 745.700 126.260 749.750 ;
        RECT 127.420 745.700 132.420 749.750 ;
        RECT 133.580 745.700 138.580 749.750 ;
        RECT 139.740 745.700 144.740 749.750 ;
        RECT 145.900 745.700 150.900 749.750 ;
        RECT 152.060 745.700 157.060 749.750 ;
        RECT 158.220 745.700 163.220 749.750 ;
        RECT 164.380 745.700 169.380 749.750 ;
        RECT 170.540 745.700 175.540 749.750 ;
        RECT 176.700 745.700 181.700 749.750 ;
        RECT 182.860 745.700 187.860 749.750 ;
        RECT 189.020 745.700 194.020 749.750 ;
        RECT 195.180 745.700 200.180 749.750 ;
        RECT 201.340 745.700 206.340 749.750 ;
        RECT 207.500 745.700 212.500 749.750 ;
        RECT 213.660 745.700 218.660 749.750 ;
        RECT 219.820 745.700 224.820 749.750 ;
        RECT 225.980 745.700 230.980 749.750 ;
        RECT 232.140 745.700 237.140 749.750 ;
        RECT 238.300 745.700 243.300 749.750 ;
        RECT 244.460 745.700 249.460 749.750 ;
        RECT 250.620 745.700 255.620 749.750 ;
        RECT 256.780 745.700 261.780 749.750 ;
        RECT 262.940 745.700 267.940 749.750 ;
        RECT 269.100 745.700 274.100 749.750 ;
        RECT 275.260 745.700 280.260 749.750 ;
        RECT 281.420 745.700 286.420 749.750 ;
        RECT 287.580 745.700 292.580 749.750 ;
        RECT 293.740 745.700 298.740 749.750 ;
        RECT 299.900 745.700 304.900 749.750 ;
        RECT 306.060 745.700 311.060 749.750 ;
        RECT 312.220 745.700 317.220 749.750 ;
        RECT 318.380 745.700 323.380 749.750 ;
        RECT 324.540 745.700 329.540 749.750 ;
        RECT 330.700 745.700 335.700 749.750 ;
        RECT 336.860 745.700 341.860 749.750 ;
        RECT 343.020 745.700 348.020 749.750 ;
        RECT 349.180 745.700 354.180 749.750 ;
        RECT 355.340 745.700 360.340 749.750 ;
        RECT 361.500 745.700 366.500 749.750 ;
        RECT 367.660 745.700 372.660 749.750 ;
        RECT 373.820 745.700 378.820 749.750 ;
        RECT 379.980 745.700 384.980 749.750 ;
        RECT 386.140 745.700 391.140 749.750 ;
        RECT 392.300 745.700 397.300 749.750 ;
        RECT 398.460 745.700 403.460 749.750 ;
        RECT 404.620 745.700 409.620 749.750 ;
        RECT 410.780 745.700 415.780 749.750 ;
        RECT 416.940 745.700 421.940 749.750 ;
        RECT 423.100 745.700 428.100 749.750 ;
        RECT 429.260 745.700 434.260 749.750 ;
        RECT 435.420 745.700 440.420 749.750 ;
        RECT 441.580 745.700 446.580 749.750 ;
        RECT 447.740 745.700 469.700 749.750 ;
        RECT 7.420 4.300 469.700 745.700 ;
        RECT 7.420 3.500 9.780 4.300 ;
        RECT 10.940 3.500 14.820 4.300 ;
        RECT 15.980 3.500 19.860 4.300 ;
        RECT 21.020 3.500 24.900 4.300 ;
        RECT 26.060 3.500 29.940 4.300 ;
        RECT 31.100 3.500 34.980 4.300 ;
        RECT 36.140 3.500 40.020 4.300 ;
        RECT 41.180 3.500 45.060 4.300 ;
        RECT 46.220 3.500 50.100 4.300 ;
        RECT 51.260 3.500 55.140 4.300 ;
        RECT 56.300 3.500 60.180 4.300 ;
        RECT 61.340 3.500 65.220 4.300 ;
        RECT 66.380 3.500 70.260 4.300 ;
        RECT 71.420 3.500 75.300 4.300 ;
        RECT 76.460 3.500 80.340 4.300 ;
        RECT 81.500 3.500 85.380 4.300 ;
        RECT 86.540 3.500 90.420 4.300 ;
        RECT 91.580 3.500 95.460 4.300 ;
        RECT 96.620 3.500 100.500 4.300 ;
        RECT 101.660 3.500 105.540 4.300 ;
        RECT 106.700 3.500 110.580 4.300 ;
        RECT 111.740 3.500 115.620 4.300 ;
        RECT 116.780 3.500 120.660 4.300 ;
        RECT 121.820 3.500 125.700 4.300 ;
        RECT 126.860 3.500 130.740 4.300 ;
        RECT 131.900 3.500 135.780 4.300 ;
        RECT 136.940 3.500 140.820 4.300 ;
        RECT 141.980 3.500 145.860 4.300 ;
        RECT 147.020 3.500 150.900 4.300 ;
        RECT 152.060 3.500 155.940 4.300 ;
        RECT 157.100 3.500 160.980 4.300 ;
        RECT 162.140 3.500 166.020 4.300 ;
        RECT 167.180 3.500 171.060 4.300 ;
        RECT 172.220 3.500 176.100 4.300 ;
        RECT 177.260 3.500 181.140 4.300 ;
        RECT 182.300 3.500 186.180 4.300 ;
        RECT 187.340 3.500 191.220 4.300 ;
        RECT 192.380 3.500 196.260 4.300 ;
        RECT 197.420 3.500 201.300 4.300 ;
        RECT 202.460 3.500 206.340 4.300 ;
        RECT 207.500 3.500 211.380 4.300 ;
        RECT 212.540 3.500 216.420 4.300 ;
        RECT 217.580 3.500 221.460 4.300 ;
        RECT 222.620 3.500 226.500 4.300 ;
        RECT 227.660 3.500 231.540 4.300 ;
        RECT 232.700 3.500 236.580 4.300 ;
        RECT 237.740 3.500 241.620 4.300 ;
        RECT 242.780 3.500 246.660 4.300 ;
        RECT 247.820 3.500 251.700 4.300 ;
        RECT 252.860 3.500 256.740 4.300 ;
        RECT 257.900 3.500 261.780 4.300 ;
        RECT 262.940 3.500 266.820 4.300 ;
        RECT 267.980 3.500 271.860 4.300 ;
        RECT 273.020 3.500 276.900 4.300 ;
        RECT 278.060 3.500 281.940 4.300 ;
        RECT 283.100 3.500 286.980 4.300 ;
        RECT 288.140 3.500 292.020 4.300 ;
        RECT 293.180 3.500 297.060 4.300 ;
        RECT 298.220 3.500 302.100 4.300 ;
        RECT 303.260 3.500 307.140 4.300 ;
        RECT 308.300 3.500 312.180 4.300 ;
        RECT 313.340 3.500 317.220 4.300 ;
        RECT 318.380 3.500 322.260 4.300 ;
        RECT 323.420 3.500 327.300 4.300 ;
        RECT 328.460 3.500 332.340 4.300 ;
        RECT 333.500 3.500 337.380 4.300 ;
        RECT 338.540 3.500 342.420 4.300 ;
        RECT 343.580 3.500 347.460 4.300 ;
        RECT 348.620 3.500 352.500 4.300 ;
        RECT 353.660 3.500 357.540 4.300 ;
        RECT 358.700 3.500 362.580 4.300 ;
        RECT 363.740 3.500 367.620 4.300 ;
        RECT 368.780 3.500 372.660 4.300 ;
        RECT 373.820 3.500 377.700 4.300 ;
        RECT 378.860 3.500 382.740 4.300 ;
        RECT 383.900 3.500 387.780 4.300 ;
        RECT 388.940 3.500 392.820 4.300 ;
        RECT 393.980 3.500 397.860 4.300 ;
        RECT 399.020 3.500 402.900 4.300 ;
        RECT 404.060 3.500 407.940 4.300 ;
        RECT 409.100 3.500 412.980 4.300 ;
        RECT 414.140 3.500 418.020 4.300 ;
        RECT 419.180 3.500 423.060 4.300 ;
        RECT 424.220 3.500 428.100 4.300 ;
        RECT 429.260 3.500 433.140 4.300 ;
        RECT 434.300 3.500 438.180 4.300 ;
        RECT 439.340 3.500 443.220 4.300 ;
        RECT 444.380 3.500 448.260 4.300 ;
        RECT 449.420 3.500 453.300 4.300 ;
        RECT 454.460 3.500 458.340 4.300 ;
        RECT 459.500 3.500 469.700 4.300 ;
      LAYER Metal3 ;
        RECT 3.500 741.740 469.190 749.700 ;
        RECT 4.300 740.580 469.190 741.740 ;
        RECT 3.500 735.580 469.190 740.580 ;
        RECT 4.300 734.420 469.190 735.580 ;
        RECT 3.500 733.900 469.190 734.420 ;
        RECT 3.500 732.740 465.700 733.900 ;
        RECT 3.500 729.420 469.190 732.740 ;
        RECT 4.300 728.260 469.190 729.420 ;
        RECT 3.500 723.260 469.190 728.260 ;
        RECT 4.300 722.700 469.190 723.260 ;
        RECT 4.300 722.100 465.700 722.700 ;
        RECT 3.500 721.540 465.700 722.100 ;
        RECT 3.500 717.100 469.190 721.540 ;
        RECT 4.300 715.940 469.190 717.100 ;
        RECT 3.500 711.500 469.190 715.940 ;
        RECT 3.500 710.940 465.700 711.500 ;
        RECT 4.300 710.340 465.700 710.940 ;
        RECT 4.300 709.780 469.190 710.340 ;
        RECT 3.500 704.780 469.190 709.780 ;
        RECT 4.300 703.620 469.190 704.780 ;
        RECT 3.500 700.300 469.190 703.620 ;
        RECT 3.500 699.140 465.700 700.300 ;
        RECT 3.500 698.620 469.190 699.140 ;
        RECT 4.300 697.460 469.190 698.620 ;
        RECT 3.500 692.460 469.190 697.460 ;
        RECT 4.300 691.300 469.190 692.460 ;
        RECT 3.500 689.100 469.190 691.300 ;
        RECT 3.500 687.940 465.700 689.100 ;
        RECT 3.500 686.300 469.190 687.940 ;
        RECT 4.300 685.140 469.190 686.300 ;
        RECT 3.500 680.140 469.190 685.140 ;
        RECT 4.300 678.980 469.190 680.140 ;
        RECT 3.500 677.900 469.190 678.980 ;
        RECT 3.500 676.740 465.700 677.900 ;
        RECT 3.500 673.980 469.190 676.740 ;
        RECT 4.300 672.820 469.190 673.980 ;
        RECT 3.500 667.820 469.190 672.820 ;
        RECT 4.300 666.700 469.190 667.820 ;
        RECT 4.300 666.660 465.700 666.700 ;
        RECT 3.500 665.540 465.700 666.660 ;
        RECT 3.500 661.660 469.190 665.540 ;
        RECT 4.300 660.500 469.190 661.660 ;
        RECT 3.500 655.500 469.190 660.500 ;
        RECT 4.300 654.340 465.700 655.500 ;
        RECT 3.500 649.340 469.190 654.340 ;
        RECT 4.300 648.180 469.190 649.340 ;
        RECT 3.500 644.300 469.190 648.180 ;
        RECT 3.500 643.180 465.700 644.300 ;
        RECT 4.300 643.140 465.700 643.180 ;
        RECT 4.300 642.020 469.190 643.140 ;
        RECT 3.500 637.020 469.190 642.020 ;
        RECT 4.300 635.860 469.190 637.020 ;
        RECT 3.500 633.100 469.190 635.860 ;
        RECT 3.500 631.940 465.700 633.100 ;
        RECT 3.500 630.860 469.190 631.940 ;
        RECT 4.300 629.700 469.190 630.860 ;
        RECT 3.500 624.700 469.190 629.700 ;
        RECT 4.300 623.540 469.190 624.700 ;
        RECT 3.500 621.900 469.190 623.540 ;
        RECT 3.500 620.740 465.700 621.900 ;
        RECT 3.500 618.540 469.190 620.740 ;
        RECT 4.300 617.380 469.190 618.540 ;
        RECT 3.500 612.380 469.190 617.380 ;
        RECT 4.300 611.220 469.190 612.380 ;
        RECT 3.500 610.700 469.190 611.220 ;
        RECT 3.500 609.540 465.700 610.700 ;
        RECT 3.500 606.220 469.190 609.540 ;
        RECT 4.300 605.060 469.190 606.220 ;
        RECT 3.500 600.060 469.190 605.060 ;
        RECT 4.300 599.500 469.190 600.060 ;
        RECT 4.300 598.900 465.700 599.500 ;
        RECT 3.500 598.340 465.700 598.900 ;
        RECT 3.500 593.900 469.190 598.340 ;
        RECT 4.300 592.740 469.190 593.900 ;
        RECT 3.500 588.300 469.190 592.740 ;
        RECT 3.500 587.740 465.700 588.300 ;
        RECT 4.300 587.140 465.700 587.740 ;
        RECT 4.300 586.580 469.190 587.140 ;
        RECT 3.500 581.580 469.190 586.580 ;
        RECT 4.300 580.420 469.190 581.580 ;
        RECT 3.500 577.100 469.190 580.420 ;
        RECT 3.500 575.940 465.700 577.100 ;
        RECT 3.500 575.420 469.190 575.940 ;
        RECT 4.300 574.260 469.190 575.420 ;
        RECT 3.500 569.260 469.190 574.260 ;
        RECT 4.300 568.100 469.190 569.260 ;
        RECT 3.500 565.900 469.190 568.100 ;
        RECT 3.500 564.740 465.700 565.900 ;
        RECT 3.500 563.100 469.190 564.740 ;
        RECT 4.300 561.940 469.190 563.100 ;
        RECT 3.500 556.940 469.190 561.940 ;
        RECT 4.300 555.780 469.190 556.940 ;
        RECT 3.500 554.700 469.190 555.780 ;
        RECT 3.500 553.540 465.700 554.700 ;
        RECT 3.500 550.780 469.190 553.540 ;
        RECT 4.300 549.620 469.190 550.780 ;
        RECT 3.500 544.620 469.190 549.620 ;
        RECT 4.300 543.500 469.190 544.620 ;
        RECT 4.300 543.460 465.700 543.500 ;
        RECT 3.500 542.340 465.700 543.460 ;
        RECT 3.500 538.460 469.190 542.340 ;
        RECT 4.300 537.300 469.190 538.460 ;
        RECT 3.500 532.300 469.190 537.300 ;
        RECT 4.300 531.140 465.700 532.300 ;
        RECT 3.500 526.140 469.190 531.140 ;
        RECT 4.300 524.980 469.190 526.140 ;
        RECT 3.500 521.100 469.190 524.980 ;
        RECT 3.500 519.980 465.700 521.100 ;
        RECT 4.300 519.940 465.700 519.980 ;
        RECT 4.300 518.820 469.190 519.940 ;
        RECT 3.500 513.820 469.190 518.820 ;
        RECT 4.300 512.660 469.190 513.820 ;
        RECT 3.500 509.900 469.190 512.660 ;
        RECT 3.500 508.740 465.700 509.900 ;
        RECT 3.500 507.660 469.190 508.740 ;
        RECT 4.300 506.500 469.190 507.660 ;
        RECT 3.500 501.500 469.190 506.500 ;
        RECT 4.300 500.340 469.190 501.500 ;
        RECT 3.500 498.700 469.190 500.340 ;
        RECT 3.500 497.540 465.700 498.700 ;
        RECT 3.500 495.340 469.190 497.540 ;
        RECT 4.300 494.180 469.190 495.340 ;
        RECT 3.500 489.180 469.190 494.180 ;
        RECT 4.300 488.020 469.190 489.180 ;
        RECT 3.500 487.500 469.190 488.020 ;
        RECT 3.500 486.340 465.700 487.500 ;
        RECT 3.500 483.020 469.190 486.340 ;
        RECT 4.300 481.860 469.190 483.020 ;
        RECT 3.500 476.860 469.190 481.860 ;
        RECT 4.300 476.300 469.190 476.860 ;
        RECT 4.300 475.700 465.700 476.300 ;
        RECT 3.500 475.140 465.700 475.700 ;
        RECT 3.500 470.700 469.190 475.140 ;
        RECT 4.300 469.540 469.190 470.700 ;
        RECT 3.500 465.100 469.190 469.540 ;
        RECT 3.500 464.540 465.700 465.100 ;
        RECT 4.300 463.940 465.700 464.540 ;
        RECT 4.300 463.380 469.190 463.940 ;
        RECT 3.500 458.380 469.190 463.380 ;
        RECT 4.300 457.220 469.190 458.380 ;
        RECT 3.500 453.900 469.190 457.220 ;
        RECT 3.500 452.740 465.700 453.900 ;
        RECT 3.500 452.220 469.190 452.740 ;
        RECT 4.300 451.060 469.190 452.220 ;
        RECT 3.500 446.060 469.190 451.060 ;
        RECT 4.300 444.900 469.190 446.060 ;
        RECT 3.500 442.700 469.190 444.900 ;
        RECT 3.500 441.540 465.700 442.700 ;
        RECT 3.500 439.900 469.190 441.540 ;
        RECT 4.300 438.740 469.190 439.900 ;
        RECT 3.500 433.740 469.190 438.740 ;
        RECT 4.300 432.580 469.190 433.740 ;
        RECT 3.500 431.500 469.190 432.580 ;
        RECT 3.500 430.340 465.700 431.500 ;
        RECT 3.500 427.580 469.190 430.340 ;
        RECT 4.300 426.420 469.190 427.580 ;
        RECT 3.500 421.420 469.190 426.420 ;
        RECT 4.300 420.300 469.190 421.420 ;
        RECT 4.300 420.260 465.700 420.300 ;
        RECT 3.500 419.140 465.700 420.260 ;
        RECT 3.500 415.260 469.190 419.140 ;
        RECT 4.300 414.100 469.190 415.260 ;
        RECT 3.500 409.100 469.190 414.100 ;
        RECT 4.300 407.940 465.700 409.100 ;
        RECT 3.500 402.940 469.190 407.940 ;
        RECT 4.300 401.780 469.190 402.940 ;
        RECT 3.500 397.900 469.190 401.780 ;
        RECT 3.500 396.780 465.700 397.900 ;
        RECT 4.300 396.740 465.700 396.780 ;
        RECT 4.300 395.620 469.190 396.740 ;
        RECT 3.500 390.620 469.190 395.620 ;
        RECT 4.300 389.460 469.190 390.620 ;
        RECT 3.500 386.700 469.190 389.460 ;
        RECT 3.500 385.540 465.700 386.700 ;
        RECT 3.500 384.460 469.190 385.540 ;
        RECT 4.300 383.300 469.190 384.460 ;
        RECT 3.500 378.300 469.190 383.300 ;
        RECT 4.300 377.140 469.190 378.300 ;
        RECT 3.500 375.500 469.190 377.140 ;
        RECT 3.500 374.340 465.700 375.500 ;
        RECT 3.500 372.140 469.190 374.340 ;
        RECT 4.300 370.980 469.190 372.140 ;
        RECT 3.500 365.980 469.190 370.980 ;
        RECT 4.300 364.820 469.190 365.980 ;
        RECT 3.500 364.300 469.190 364.820 ;
        RECT 3.500 363.140 465.700 364.300 ;
        RECT 3.500 359.820 469.190 363.140 ;
        RECT 4.300 358.660 469.190 359.820 ;
        RECT 3.500 353.660 469.190 358.660 ;
        RECT 4.300 353.100 469.190 353.660 ;
        RECT 4.300 352.500 465.700 353.100 ;
        RECT 3.500 351.940 465.700 352.500 ;
        RECT 3.500 347.500 469.190 351.940 ;
        RECT 4.300 346.340 469.190 347.500 ;
        RECT 3.500 341.900 469.190 346.340 ;
        RECT 3.500 341.340 465.700 341.900 ;
        RECT 4.300 340.740 465.700 341.340 ;
        RECT 4.300 340.180 469.190 340.740 ;
        RECT 3.500 335.180 469.190 340.180 ;
        RECT 4.300 334.020 469.190 335.180 ;
        RECT 3.500 330.700 469.190 334.020 ;
        RECT 3.500 329.540 465.700 330.700 ;
        RECT 3.500 329.020 469.190 329.540 ;
        RECT 4.300 327.860 469.190 329.020 ;
        RECT 3.500 322.860 469.190 327.860 ;
        RECT 4.300 321.700 469.190 322.860 ;
        RECT 3.500 319.500 469.190 321.700 ;
        RECT 3.500 318.340 465.700 319.500 ;
        RECT 3.500 316.700 469.190 318.340 ;
        RECT 4.300 315.540 469.190 316.700 ;
        RECT 3.500 310.540 469.190 315.540 ;
        RECT 4.300 309.380 469.190 310.540 ;
        RECT 3.500 308.300 469.190 309.380 ;
        RECT 3.500 307.140 465.700 308.300 ;
        RECT 3.500 304.380 469.190 307.140 ;
        RECT 4.300 303.220 469.190 304.380 ;
        RECT 3.500 298.220 469.190 303.220 ;
        RECT 4.300 297.100 469.190 298.220 ;
        RECT 4.300 297.060 465.700 297.100 ;
        RECT 3.500 295.940 465.700 297.060 ;
        RECT 3.500 292.060 469.190 295.940 ;
        RECT 4.300 290.900 469.190 292.060 ;
        RECT 3.500 285.900 469.190 290.900 ;
        RECT 4.300 284.740 465.700 285.900 ;
        RECT 3.500 279.740 469.190 284.740 ;
        RECT 4.300 278.580 469.190 279.740 ;
        RECT 3.500 274.700 469.190 278.580 ;
        RECT 3.500 273.580 465.700 274.700 ;
        RECT 4.300 273.540 465.700 273.580 ;
        RECT 4.300 272.420 469.190 273.540 ;
        RECT 3.500 267.420 469.190 272.420 ;
        RECT 4.300 266.260 469.190 267.420 ;
        RECT 3.500 263.500 469.190 266.260 ;
        RECT 3.500 262.340 465.700 263.500 ;
        RECT 3.500 261.260 469.190 262.340 ;
        RECT 4.300 260.100 469.190 261.260 ;
        RECT 3.500 255.100 469.190 260.100 ;
        RECT 4.300 253.940 469.190 255.100 ;
        RECT 3.500 252.300 469.190 253.940 ;
        RECT 3.500 251.140 465.700 252.300 ;
        RECT 3.500 248.940 469.190 251.140 ;
        RECT 4.300 247.780 469.190 248.940 ;
        RECT 3.500 242.780 469.190 247.780 ;
        RECT 4.300 241.620 469.190 242.780 ;
        RECT 3.500 241.100 469.190 241.620 ;
        RECT 3.500 239.940 465.700 241.100 ;
        RECT 3.500 236.620 469.190 239.940 ;
        RECT 4.300 235.460 469.190 236.620 ;
        RECT 3.500 230.460 469.190 235.460 ;
        RECT 4.300 229.900 469.190 230.460 ;
        RECT 4.300 229.300 465.700 229.900 ;
        RECT 3.500 228.740 465.700 229.300 ;
        RECT 3.500 224.300 469.190 228.740 ;
        RECT 4.300 223.140 469.190 224.300 ;
        RECT 3.500 218.700 469.190 223.140 ;
        RECT 3.500 218.140 465.700 218.700 ;
        RECT 4.300 217.540 465.700 218.140 ;
        RECT 4.300 216.980 469.190 217.540 ;
        RECT 3.500 211.980 469.190 216.980 ;
        RECT 4.300 210.820 469.190 211.980 ;
        RECT 3.500 207.500 469.190 210.820 ;
        RECT 3.500 206.340 465.700 207.500 ;
        RECT 3.500 205.820 469.190 206.340 ;
        RECT 4.300 204.660 469.190 205.820 ;
        RECT 3.500 199.660 469.190 204.660 ;
        RECT 4.300 198.500 469.190 199.660 ;
        RECT 3.500 196.300 469.190 198.500 ;
        RECT 3.500 195.140 465.700 196.300 ;
        RECT 3.500 193.500 469.190 195.140 ;
        RECT 4.300 192.340 469.190 193.500 ;
        RECT 3.500 187.340 469.190 192.340 ;
        RECT 4.300 186.180 469.190 187.340 ;
        RECT 3.500 185.100 469.190 186.180 ;
        RECT 3.500 183.940 465.700 185.100 ;
        RECT 3.500 181.180 469.190 183.940 ;
        RECT 4.300 180.020 469.190 181.180 ;
        RECT 3.500 175.020 469.190 180.020 ;
        RECT 4.300 173.900 469.190 175.020 ;
        RECT 4.300 173.860 465.700 173.900 ;
        RECT 3.500 172.740 465.700 173.860 ;
        RECT 3.500 168.860 469.190 172.740 ;
        RECT 4.300 167.700 469.190 168.860 ;
        RECT 3.500 162.700 469.190 167.700 ;
        RECT 4.300 161.540 465.700 162.700 ;
        RECT 3.500 156.540 469.190 161.540 ;
        RECT 4.300 155.380 469.190 156.540 ;
        RECT 3.500 151.500 469.190 155.380 ;
        RECT 3.500 150.380 465.700 151.500 ;
        RECT 4.300 150.340 465.700 150.380 ;
        RECT 4.300 149.220 469.190 150.340 ;
        RECT 3.500 144.220 469.190 149.220 ;
        RECT 4.300 143.060 469.190 144.220 ;
        RECT 3.500 140.300 469.190 143.060 ;
        RECT 3.500 139.140 465.700 140.300 ;
        RECT 3.500 138.060 469.190 139.140 ;
        RECT 4.300 136.900 469.190 138.060 ;
        RECT 3.500 131.900 469.190 136.900 ;
        RECT 4.300 130.740 469.190 131.900 ;
        RECT 3.500 129.100 469.190 130.740 ;
        RECT 3.500 127.940 465.700 129.100 ;
        RECT 3.500 125.740 469.190 127.940 ;
        RECT 4.300 124.580 469.190 125.740 ;
        RECT 3.500 119.580 469.190 124.580 ;
        RECT 4.300 118.420 469.190 119.580 ;
        RECT 3.500 117.900 469.190 118.420 ;
        RECT 3.500 116.740 465.700 117.900 ;
        RECT 3.500 113.420 469.190 116.740 ;
        RECT 4.300 112.260 469.190 113.420 ;
        RECT 3.500 107.260 469.190 112.260 ;
        RECT 4.300 106.700 469.190 107.260 ;
        RECT 4.300 106.100 465.700 106.700 ;
        RECT 3.500 105.540 465.700 106.100 ;
        RECT 3.500 101.100 469.190 105.540 ;
        RECT 4.300 99.940 469.190 101.100 ;
        RECT 3.500 95.500 469.190 99.940 ;
        RECT 3.500 94.940 465.700 95.500 ;
        RECT 4.300 94.340 465.700 94.940 ;
        RECT 4.300 93.780 469.190 94.340 ;
        RECT 3.500 88.780 469.190 93.780 ;
        RECT 4.300 87.620 469.190 88.780 ;
        RECT 3.500 84.300 469.190 87.620 ;
        RECT 3.500 83.140 465.700 84.300 ;
        RECT 3.500 82.620 469.190 83.140 ;
        RECT 4.300 81.460 469.190 82.620 ;
        RECT 3.500 76.460 469.190 81.460 ;
        RECT 4.300 75.300 469.190 76.460 ;
        RECT 3.500 73.100 469.190 75.300 ;
        RECT 3.500 71.940 465.700 73.100 ;
        RECT 3.500 70.300 469.190 71.940 ;
        RECT 4.300 69.140 469.190 70.300 ;
        RECT 3.500 64.140 469.190 69.140 ;
        RECT 4.300 62.980 469.190 64.140 ;
        RECT 3.500 61.900 469.190 62.980 ;
        RECT 3.500 60.740 465.700 61.900 ;
        RECT 3.500 57.980 469.190 60.740 ;
        RECT 4.300 56.820 469.190 57.980 ;
        RECT 3.500 51.820 469.190 56.820 ;
        RECT 4.300 50.700 469.190 51.820 ;
        RECT 4.300 50.660 465.700 50.700 ;
        RECT 3.500 49.540 465.700 50.660 ;
        RECT 3.500 45.660 469.190 49.540 ;
        RECT 4.300 44.500 469.190 45.660 ;
        RECT 3.500 39.500 469.190 44.500 ;
        RECT 4.300 38.340 465.700 39.500 ;
        RECT 3.500 33.340 469.190 38.340 ;
        RECT 4.300 32.180 469.190 33.340 ;
        RECT 3.500 28.300 469.190 32.180 ;
        RECT 3.500 27.180 465.700 28.300 ;
        RECT 4.300 27.140 465.700 27.180 ;
        RECT 4.300 26.020 469.190 27.140 ;
        RECT 3.500 21.020 469.190 26.020 ;
        RECT 4.300 19.860 469.190 21.020 ;
        RECT 3.500 17.100 469.190 19.860 ;
        RECT 3.500 15.940 465.700 17.100 ;
        RECT 3.500 14.860 469.190 15.940 ;
        RECT 4.300 13.700 469.190 14.860 ;
        RECT 3.500 8.700 469.190 13.700 ;
        RECT 4.300 7.980 469.190 8.700 ;
      LAYER Metal4 ;
        RECT 5.180 733.640 462.980 746.390 ;
        RECT 5.180 16.890 21.940 733.640 ;
        RECT 24.140 16.890 25.240 733.640 ;
        RECT 27.440 16.890 98.740 733.640 ;
        RECT 100.940 16.890 102.040 733.640 ;
        RECT 104.240 16.890 175.540 733.640 ;
        RECT 177.740 16.890 178.840 733.640 ;
        RECT 181.040 16.890 252.340 733.640 ;
        RECT 254.540 16.890 255.640 733.640 ;
        RECT 257.840 16.890 329.140 733.640 ;
        RECT 331.340 16.890 332.440 733.640 ;
        RECT 334.640 16.890 405.940 733.640 ;
        RECT 408.140 16.890 409.240 733.640 ;
        RECT 411.440 16.890 462.980 733.640 ;
      LAYER Metal5 ;
        RECT 5.100 698.090 463.060 739.700 ;
        RECT 5.100 695.490 5.920 698.090 ;
        RECT 5.100 658.990 463.060 695.490 ;
        RECT 5.100 656.390 5.920 658.990 ;
        RECT 5.100 619.890 463.060 656.390 ;
        RECT 5.100 617.290 5.920 619.890 ;
        RECT 5.100 580.790 463.060 617.290 ;
        RECT 5.100 578.190 5.920 580.790 ;
        RECT 5.100 541.690 463.060 578.190 ;
        RECT 5.100 539.090 5.920 541.690 ;
        RECT 5.100 502.590 463.060 539.090 ;
        RECT 5.100 499.990 5.920 502.590 ;
        RECT 5.100 463.490 463.060 499.990 ;
        RECT 5.100 460.890 5.920 463.490 ;
        RECT 5.100 424.390 463.060 460.890 ;
        RECT 5.100 421.790 5.920 424.390 ;
        RECT 5.100 385.290 463.060 421.790 ;
        RECT 5.100 382.690 5.920 385.290 ;
        RECT 5.100 346.190 463.060 382.690 ;
        RECT 5.100 343.590 5.920 346.190 ;
        RECT 5.100 307.090 463.060 343.590 ;
        RECT 5.100 304.490 5.920 307.090 ;
        RECT 5.100 267.990 463.060 304.490 ;
        RECT 5.100 265.390 5.920 267.990 ;
        RECT 5.100 228.890 463.060 265.390 ;
        RECT 5.100 226.290 5.920 228.890 ;
        RECT 5.100 189.790 463.060 226.290 ;
        RECT 5.100 187.190 5.920 189.790 ;
        RECT 5.100 150.690 463.060 187.190 ;
        RECT 5.100 148.090 5.920 150.690 ;
        RECT 5.100 111.590 463.060 148.090 ;
        RECT 5.100 108.990 5.920 111.590 ;
        RECT 5.100 72.490 463.060 108.990 ;
        RECT 5.100 69.890 5.920 72.490 ;
        RECT 5.100 33.390 463.060 69.890 ;
        RECT 5.100 30.790 5.920 33.390 ;
        RECT 5.100 16.860 463.060 30.790 ;
  END
END housekeeping
END LIBRARY

