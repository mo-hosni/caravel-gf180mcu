* NGSPICE file created from mprj_io_buffer.ext - technology: gf180mcuC

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__fill_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__fill_1 VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__fill_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__fill_2 VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__clkbuf_8 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__clkbuf_8 I Z VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__fillcap_4 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__fillcap_4 VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__antenna abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__antenna I VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__fillcap_8 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__fillcap_8 VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__endcap abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__endcap VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__fillcap_32 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__fillcap_32 VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__fillcap_16 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__fillcap_16 VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__filltie abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__filltie VDD VSS
.ends

.subckt mprj_io_buffer VDD VSS mgmt_gpio_in[0] mgmt_gpio_in[10] mgmt_gpio_in[11] mgmt_gpio_in[12]
+ mgmt_gpio_in[13] mgmt_gpio_in[14] mgmt_gpio_in[15] mgmt_gpio_in[16] mgmt_gpio_in[17]
+ mgmt_gpio_in[1] mgmt_gpio_in[2] mgmt_gpio_in[3] mgmt_gpio_in[4] mgmt_gpio_in[5]
+ mgmt_gpio_in[6] mgmt_gpio_in[7] mgmt_gpio_in[8] mgmt_gpio_in[9] mgmt_gpio_in_buf[0]
+ mgmt_gpio_in_buf[10] mgmt_gpio_in_buf[11] mgmt_gpio_in_buf[12] mgmt_gpio_in_buf[13]
+ mgmt_gpio_in_buf[14] mgmt_gpio_in_buf[15] mgmt_gpio_in_buf[16] mgmt_gpio_in_buf[17]
+ mgmt_gpio_in_buf[1] mgmt_gpio_in_buf[2] mgmt_gpio_in_buf[3] mgmt_gpio_in_buf[4]
+ mgmt_gpio_in_buf[5] mgmt_gpio_in_buf[6] mgmt_gpio_in_buf[7] mgmt_gpio_in_buf[8]
+ mgmt_gpio_in_buf[9] mgmt_gpio_oeb[0] mgmt_gpio_oeb[1] mgmt_gpio_oeb_buf[0] mgmt_gpio_oeb_buf[1]
+ mgmt_gpio_out[0] mgmt_gpio_out[10] mgmt_gpio_out[11] mgmt_gpio_out[12] mgmt_gpio_out[13]
+ mgmt_gpio_out[14] mgmt_gpio_out[15] mgmt_gpio_out[16] mgmt_gpio_out[17] mgmt_gpio_out[1]
+ mgmt_gpio_out[2] mgmt_gpio_out[3] mgmt_gpio_out[4] mgmt_gpio_out[5] mgmt_gpio_out[6]
+ mgmt_gpio_out[7] mgmt_gpio_out[8] mgmt_gpio_out[9] mgmt_gpio_out_buf[0] mgmt_gpio_out_buf[10]
+ mgmt_gpio_out_buf[11] mgmt_gpio_out_buf[12] mgmt_gpio_out_buf[13] mgmt_gpio_out_buf[14]
+ mgmt_gpio_out_buf[15] mgmt_gpio_out_buf[16] mgmt_gpio_out_buf[17] mgmt_gpio_out_buf[1]
+ mgmt_gpio_out_buf[2] mgmt_gpio_out_buf[3] mgmt_gpio_out_buf[4] mgmt_gpio_out_buf[5]
+ mgmt_gpio_out_buf[6] mgmt_gpio_out_buf[7] mgmt_gpio_out_buf[8] mgmt_gpio_out_buf[9]
XFILLER_3_67 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_9_77 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XBUF\[28\] mgmt_gpio_in[8] mgmt_gpio_in_buf[8] VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_8
XBUF\[5\] mgmt_gpio_out[5] mgmt_gpio_out_buf[5] VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_8
XFILLER_2_143 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_6_56 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_6_34 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_9_138 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XBUF\[10\] mgmt_gpio_out[10] mgmt_gpio_out_buf[10] VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_8
XFILLER_3_57 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_10_104 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_6_108 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_5_141 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_9_12 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_69 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_3_2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_BUF\[19\]_I mgmt_gpio_oeb[1] VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_BUF\[37\]_I mgmt_gpio_in[17] VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_BUF\[28\]_I mgmt_gpio_in[8] VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_10_138 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_9_106 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_BUF\[4\]_I mgmt_gpio_out[4] VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_9_79 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_5_131 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_37 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_2_101 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XBUF\[33\] mgmt_gpio_in[13] mgmt_gpio_in_buf[13] VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_8
XBUF\[3\] mgmt_gpio_out[3] mgmt_gpio_out_buf[3] VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_8
XBUF\[26\] mgmt_gpio_in[6] mgmt_gpio_in_buf[6] VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_8
XFILLER_2_135 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_6_37 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_6_48 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_1_70 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_10_107 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_5_144 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XBUF\[19\] mgmt_gpio_oeb[1] mgmt_gpio_oeb_buf[1] VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_8
XFILLER_1_2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA_BUF\[7\]_I mgmt_gpio_out[7] VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XBUF\[31\] mgmt_gpio_in[11] mgmt_gpio_in_buf[11] VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_8
XFILLER_8_143 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_7_93 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_0 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_3_29 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_9_39 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_2_105 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XBUF\[24\] mgmt_gpio_in[4] mgmt_gpio_in_buf[4] VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_8
XFILLER_1_73 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_1_84 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XBUF\[1\] mgmt_gpio_out[1] mgmt_gpio_out_buf[1] VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_8
XFILLER_7_61 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_8_100 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_BUF\[30\]_I mgmt_gpio_in[10] VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_5_103 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_BUF\[12\]_I mgmt_gpio_out[12] VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_BUF\[21\]_I mgmt_gpio_in[1] VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_4_40 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_2_139 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_10_72 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_10_61 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XBUF\[17\] mgmt_gpio_out[17] mgmt_gpio_out_buf[17] VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_8
XFILLER_7_95 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_7_73 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XPHY_2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_1_42 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_8_135 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_8_102 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_4_42 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_1_141 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_2_108 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_10_41 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_1_10 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_1_76 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XBUF\[22\] mgmt_gpio_in[2] mgmt_gpio_in_buf[2] VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_8
XANTENNA_BUF\[24\]_I mgmt_gpio_in[4] VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_BUF\[33\]_I mgmt_gpio_in[13] VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_4 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA_BUF\[15\]_I mgmt_gpio_out[15] VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_5_139 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_BUF\[0\]_I mgmt_gpio_out[0] VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XBUF\[15\] mgmt_gpio_out[15] mgmt_gpio_out_buf[15] VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_8
XFILLER_7_65 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_5 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_8_2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_4_99 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_7_33 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_6 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_8_105 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_4_34 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_1_111 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_1_144 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_BUF\[36\]_I mgmt_gpio_in[16] VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_BUF\[18\]_I mgmt_gpio_oeb[0] VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_BUF\[27\]_I mgmt_gpio_in[7] VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_8_139 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_7_89 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_7 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XBUF\[20\] mgmt_gpio_in[0] mgmt_gpio_in_buf[0] VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_8
XANTENNA_BUF\[3\]_I mgmt_gpio_out[3] VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_10_45 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_10_34 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XBUF\[8\] mgmt_gpio_out[8] mgmt_gpio_out_buf[8] VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_8
XFILLER_1_14 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_8 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XBUF\[13\] mgmt_gpio_out[13] mgmt_gpio_out_buf[13] VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_8
XFILLER_4_143 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_4_69 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_6_2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_8_108 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_7_69 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_9 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_8_6 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_4_37 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_10_69 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XBUF\[36\] mgmt_gpio_in[16] mgmt_gpio_in_buf[16] VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_8
XANTENNA_BUF\[6\]_I mgmt_gpio_out[6] VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_5_70 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_10_37 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XBUF\[6\] mgmt_gpio_out[6] mgmt_gpio_out_buf[6] VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_8
XBUF\[29\] mgmt_gpio_in[9] mgmt_gpio_in_buf[9] VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_8
XFILLER_4_135 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XBUF\[11\] mgmt_gpio_out[11] mgmt_gpio_out_buf[11] VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_8
XTAP_40 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_4_2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_7_144 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_7_122 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_BUF\[20\]_I mgmt_gpio_in[0] VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_BUF\[11\]_I mgmt_gpio_out[11] VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_1_139 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_41 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_6_6 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_30 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA_BUF\[9\]_I mgmt_gpio_out[9] VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XBUF\[34\] mgmt_gpio_in[14] mgmt_gpio_in_buf[14] VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_8
XFILLER_2_40 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_5_73 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_42 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_31 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XBUF\[4\] mgmt_gpio_out[4] mgmt_gpio_out_buf[4] VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_8
XFILLER_2_96 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XBUF\[27\] mgmt_gpio_in[7] mgmt_gpio_in_buf[7] VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_8
XFILLER_8_40 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_8_84 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_4_105 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_43 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_32 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA_BUF\[14\]_I mgmt_gpio_out[14] VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_BUF\[23\]_I mgmt_gpio_in[3] VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_2_2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_BUF\[32\]_I mgmt_gpio_in[12] VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_8_96 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_8_52 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_4_139 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_5_42 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_142 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_44 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_33 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_4_6 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_22 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_2_98 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_7_126 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XBUF\[32\] mgmt_gpio_in[12] mgmt_gpio_in_buf[12] VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_8
XTAP_45 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_10_2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_34 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_5_10 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_23 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XBUF\[2\] mgmt_gpio_out[2] mgmt_gpio_out_buf[2] VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_8
XBUF\[25\] mgmt_gpio_in[5] mgmt_gpio_in_buf[5] VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_8
XFILLER_4_108 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_144 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_46 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA_BUF\[26\]_I mgmt_gpio_in[6] VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_35 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA_BUF\[35\]_I mgmt_gpio_in[15] VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_24 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_2_34 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_BUF\[17\]_I mgmt_gpio_out[17] VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XBUF\[18\] mgmt_gpio_oeb[0] mgmt_gpio_oeb_buf[0] VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_8
XFILLER_8_88 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_8_44 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_BUF\[2\]_I mgmt_gpio_out[2] VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_47 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_36 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_134 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_25 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_20 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_2_6 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_2_68 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_8_56 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_8_34 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XBUF\[30\] mgmt_gpio_in[10] mgmt_gpio_in_buf[10] VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_8
XPHY_21 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_37 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_10 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_26 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XBUF\[23\] mgmt_gpio_in[3] mgmt_gpio_in_buf[3] VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_8
XFILLER_3_144 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_3_122 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XBUF\[0\] mgmt_gpio_out[0] mgmt_gpio_out_buf[0] VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_8
XFILLER_10_6 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_38 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_5_14 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_103 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_27 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_11 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_2_37 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_BUF\[29\]_I mgmt_gpio_in[9] VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_BUF\[5\]_I mgmt_gpio_out[5] VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_3_80 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XBUF\[16\] mgmt_gpio_out[16] mgmt_gpio_out_buf[16] VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_8
XTAP_39 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_12 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_28 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_9_2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_8_37 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_6_143 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_6 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_3_70 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_138 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_13 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_6_92 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_29 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_6_100 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_9_70 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_BUF\[10\]_I mgmt_gpio_out[10] VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XBUF\[21\] mgmt_gpio_in[1] mgmt_gpio_in_buf[1] VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_8
XFILLER_0_72 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_6_60 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XBUF\[9\] mgmt_gpio_out[9] mgmt_gpio_out_buf[9] VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_8
XANTENNA_BUF\[8\]_I mgmt_gpio_out[8] VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_14 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_3_126 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_3_61 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XBUF\[14\] mgmt_gpio_out[14] mgmt_gpio_out_buf[14] VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_8
XFILLER_0_107 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_15 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_7_2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_3_73 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_10_142 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_6_135 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_6_102 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_BUF\[22\]_I mgmt_gpio_in[2] VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_16 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_6_40 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_BUF\[31\]_I mgmt_gpio_in[11] VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_9_144 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_BUF\[13\]_I mgmt_gpio_out[13] VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XBUF\[37\] mgmt_gpio_in[17] mgmt_gpio_in_buf[17] VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_8
XFILLER_9_73 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_17 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_9_134 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XBUF\[7\] mgmt_gpio_out[7] mgmt_gpio_out_buf[7] VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_8
XFILLER_10_144 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_3_118 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_65 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XBUF\[12\] mgmt_gpio_out[12] mgmt_gpio_out_buf[12] VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_8
XPHY_18 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_10_134 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_6_105 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_5_2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_3_65 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_3_76 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_99 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_19 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA_BUF\[34\]_I mgmt_gpio_in[14] VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_BUF\[25\]_I mgmt_gpio_in[5] VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_7_6 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_3_88 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA_BUF\[16\]_I mgmt_gpio_out[16] VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_6_139 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XBUF\[35\] mgmt_gpio_in[15] mgmt_gpio_in_buf[15] VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_8
XANTENNA_BUF\[1\]_I mgmt_gpio_out[1] VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_9_43 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_9_10 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_34 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_6_88 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_6_44 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
.ends

